* NGSPICE file created from r2r_dac_control.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VPWR VGND 0.545943f
C1 VPB VGND 0.116247f
C2 VPWR VPB 0.078686f
C3 VPWR VNB 0.61942f
C4 VGND VNB 0.553666f
C5 VPB VNB 0.427572f
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
C0 VPB VGND 0.349732f
C1 VPB VPWR 0.136888f
C2 VPWR VGND 1.56539f
C3 VPWR VNB 1.67352f
C4 VGND VNB 1.46552f
C5 VPB VNB 1.13634f
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
C0 VPB VGND 0.219503f
C1 VPB VPWR 0.104823f
C2 VPWR VGND 1.27274f
C3 VPWR VNB 1.14152f
C4 VGND VNB 0.991595f
C5 VPB VNB 0.781956f
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
C0 VPB VGND 0.079664f
C1 VPB VPWR 0.062496f
C2 VPWR VGND 0.352999f
C3 VPWR VNB 0.469966f
C4 VGND VNB 0.427318f
C5 VPB VNB 0.338976f
.ends

.subckt sky130_fd_sc_hd__dfxtp_4 VGND VPWR VNB VPB Q D CLK a_1020_47# a_975_413# a_891_413#
+ a_193_47# a_381_47# a_1062_300# a_572_47# a_568_413# a_475_413# a_634_183# a_27_47#
X0 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X1 a_1020_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X2 a_572_47# a_193_47# a_475_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X3 VPWR a_1062_300# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.09135 ps=0.855 w=0.42 l=0.15
X4 a_634_183# a_475_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X5 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_475_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8 VGND a_1062_300# a_1020_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X9 VPWR a_634_183# a_568_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X11 a_568_413# a_27_47# a_475_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X12 a_634_183# a_475_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_183# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X17 VGND a_891_413# a_1062_300# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X18 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 VPWR a_891_413# a_1062_300# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.28 ps=2.56 w=1 l=0.15
X25 a_891_413# a_193_47# a_634_183# VNB sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X26 a_475_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X27 VGND a_634_183# a_572_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
C0 a_1020_47# VPWR 4.79e-19
C1 a_1020_47# VGND 0.004151f
C2 a_1062_300# a_1020_47# 8.75e-20
C3 a_572_47# a_193_47# 0.001131f
C4 a_975_413# VPWR 0.00475f
C5 a_193_47# a_27_47# 0.723863f
C6 VPB a_193_47# 0.141384f
C7 a_572_47# a_634_183# 6.29e-20
C8 a_1020_47# a_891_413# 0.00605f
C9 VGND a_975_413# 5.62e-19
C10 a_634_183# a_27_47# 0.166122f
C11 VPB a_634_183# 0.073615f
C12 a_568_413# VPWR 0.002673f
C13 CLK a_27_47# 0.21376f
C14 VPB CLK 0.070057f
C15 a_568_413# a_475_413# 0.007015f
C16 a_381_47# a_568_413# 0.001089f
C17 a_975_413# a_891_413# 0.008802f
C18 VPWR a_27_47# 0.383097f
C19 VGND a_572_47# 0.003976f
C20 VPB VPWR 0.198564f
C21 a_572_47# a_475_413# 0.006375f
C22 VGND a_27_47# 0.12468f
C23 a_475_413# a_27_47# 0.178436f
C24 a_193_47# a_634_183# 0.130991f
C25 VGND VPB 0.014659f
C26 a_381_47# a_572_47# 1.46e-19
C27 VPB a_475_413# 0.075941f
C28 D a_27_47# 0.096989f
C29 Q a_27_47# 3.44e-19
C30 VPB D 0.09609f
C31 a_381_47# a_27_47# 0.03397f
C32 Q VPB 0.013356f
C33 a_381_47# VPB 0.013583f
C34 a_1062_300# a_27_47# 0.048687f
C35 a_193_47# CLK 0.001315f
C36 a_1062_300# VPB 0.24732f
C37 a_891_413# a_27_47# 0.037767f
C38 a_891_413# VPB 0.068757f
C39 a_193_47# VPWR 0.106627f
C40 VGND a_193_47# 0.305428f
C41 VPWR a_634_183# 0.102093f
C42 a_193_47# a_475_413# 0.157543f
C43 a_193_47# D 0.103962f
C44 Q a_193_47# 4.61e-19
C45 VGND a_634_183# 0.123913f
C46 a_381_47# a_193_47# 0.16187f
C47 a_475_413# a_634_183# 0.248641f
C48 a_1062_300# a_193_47# 0.030243f
C49 VPWR CLK 0.019411f
C50 a_381_47# a_634_183# 3.45e-19
C51 VGND CLK 0.019463f
C52 a_1062_300# a_634_183# 1.25e-19
C53 a_891_413# a_193_47# 0.139283f
C54 a_891_413# a_634_183# 0.035483f
C55 VGND VPWR 0.100633f
C56 VPWR a_475_413# 0.168224f
C57 VPWR D 0.027256f
C58 Q VPWR 0.335782f
C59 a_381_47# VPWR 0.053383f
C60 VGND a_475_413# 0.09216f
C61 VGND D 0.026396f
C62 VGND Q 0.242058f
C63 a_568_413# a_27_47# 0.002418f
C64 a_1062_300# VPWR 0.226048f
C65 a_381_47# VGND 0.044834f
C66 a_381_47# a_475_413# 0.035644f
C67 a_1020_47# a_634_183# 3.37e-20
C68 a_1062_300# VGND 0.194826f
C69 a_381_47# D 0.076792f
C70 a_1062_300# Q 0.387919f
C71 a_891_413# VPWR 0.113945f
C72 VGND a_891_413# 0.116731f
C73 a_572_47# a_27_47# 7.78e-20
C74 a_975_413# a_193_47# 2.81e-19
C75 a_891_413# Q 0.001398f
C76 VPB a_27_47# 0.275432f
C77 a_975_413# a_634_183# 9.88e-19
C78 a_1062_300# a_891_413# 0.285494f
C79 Q VNB 0.060797f
C80 VGND VNB 0.988933f
C81 VPWR VNB 0.823111f
C82 D VNB 0.129726f
C83 CLK VNB 0.195983f
C84 VPB VNB 1.75651f
C85 a_381_47# VNB 0.016397f
C86 a_891_413# VNB 0.160892f
C87 a_1062_300# VNB 0.529662f
C88 a_475_413# VNB 0.137184f
C89 a_634_183# VNB 0.150209f
C90 a_193_47# VNB 0.271178f
C91 a_27_47# VNB 0.468295f
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VNB VPB VGND VPWR A X a_110_47#
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
C0 VPB a_110_47# 0.527557f
C1 VPWR a_110_47# 0.669976f
C2 X a_110_47# 1.62234f
C3 A a_110_47# 0.306578f
C4 VGND a_110_47# 0.512392f
C5 VPWR VPB 0.183858f
C6 X VPB 0.03148f
C7 VPB A 0.133397f
C8 VGND VPB 0.011388f
C9 X VPWR 1.36494f
C10 VPWR A 0.111641f
C11 VGND VPWR 0.187357f
C12 X A 0.002918f
C13 X VGND 0.976879f
C14 VGND A 0.115353f
C15 VGND VNB 1.01442f
C16 X VNB 0.110579f
C17 VPWR VNB 0.834786f
C18 A VNB 0.494734f
C19 VPB VNB 1.84511f
C20 a_110_47# VNB 1.73295f
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR VPB VNB CLK D RESET_B Q a_1462_47# a_543_47#
+ a_651_413# a_193_47# a_805_47# a_448_47# a_639_47# a_1283_21# a_761_289# a_1108_47#
+ a_1217_47# a_1270_413# a_27_47#
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
C0 a_805_47# RESET_B 0.003155f
C1 a_651_413# a_543_47# 0.057222f
C2 CLK VPWR 0.017406f
C3 VPWR Q 0.099692f
C4 VPB CLK 0.069345f
C5 VPB Q 0.011004f
C6 CLK a_27_47# 0.233602f
C7 a_651_413# RESET_B 0.012196f
C8 a_193_47# CLK 7.94e-19
C9 Q a_27_47# 2.63e-20
C10 a_1462_47# VGND 0.002215f
C11 a_193_47# Q 1.81e-19
C12 VPWR a_761_289# 0.10497f
C13 VPB a_761_289# 0.099418f
C14 a_1462_47# a_1283_21# 0.007399f
C15 a_761_289# a_27_47# 0.07009f
C16 a_193_47# a_761_289# 0.186387f
C17 VPWR VGND 0.050202f
C18 VPB VGND 0.009994f
C19 a_1283_21# VPWR 0.208909f
C20 VGND a_27_47# 0.253961f
C21 VGND D 0.051614f
C22 a_193_47# VGND 0.063057f
C23 a_1108_47# VPWR 0.17338f
C24 VPB a_1283_21# 0.136539f
C25 VPWR a_1270_413# 7.19e-19
C26 VPWR a_543_47# 0.100285f
C27 a_448_47# VPWR 0.068142f
C28 a_1283_21# a_27_47# 0.043567f
C29 a_1108_47# VPB 0.113409f
C30 a_193_47# a_1283_21# 0.042415f
C31 a_1462_47# RESET_B 0.002879f
C32 a_1108_47# a_27_47# 0.102355f
C33 VPB a_543_47# 0.095793f
C34 a_448_47# VPB 0.014137f
C35 a_1108_47# a_193_47# 0.125324f
C36 a_193_47# a_1270_413# 1.46e-19
C37 a_543_47# a_27_47# 0.115353f
C38 a_543_47# D 7.35e-20
C39 a_448_47# a_27_47# 0.093133f
C40 a_448_47# D 0.155634f
C41 a_193_47# a_543_47# 0.229804f
C42 a_1217_47# a_27_47# 2.56e-19
C43 a_448_47# a_193_47# 0.064178f
C44 a_1217_47# a_193_47# 2.36e-20
C45 a_639_47# a_27_47# 0.001881f
C46 VPWR RESET_B 0.065186f
C47 a_639_47# a_193_47# 2.28e-19
C48 VPB RESET_B 0.138482f
C49 a_27_47# RESET_B 0.296336f
C50 RESET_B D 4.72e-19
C51 CLK VGND 0.017208f
C52 a_193_47# RESET_B 0.026903f
C53 VGND Q 0.061585f
C54 a_651_413# VPWR 0.12856f
C55 a_1283_21# Q 0.059778f
C56 a_761_289# VGND 0.073384f
C57 a_651_413# VPB 0.013543f
C58 a_1108_47# Q 9.8e-19
C59 a_651_413# a_27_47# 9.73e-19
C60 a_651_413# a_193_47# 0.034619f
C61 a_1108_47# a_761_289# 0.051162f
C62 a_761_289# a_1270_413# 2.6e-19
C63 a_761_289# a_543_47# 0.209641f
C64 a_1217_47# a_761_289# 4.2e-19
C65 CLK RESET_B 1.09e-19
C66 a_1283_21# VGND 0.239533f
C67 Q RESET_B 9.12e-19
C68 a_639_47# a_761_289# 3.16e-19
C69 a_1108_47# VGND 0.148001f
C70 VGND a_543_47# 0.122935f
C71 a_448_47# VGND 0.0661f
C72 a_1217_47# VGND 9.68e-19
C73 a_1108_47# a_1283_21# 0.233657f
C74 a_761_289# RESET_B 0.166114f
C75 a_639_47# VGND 0.008634f
C76 a_805_47# a_761_289# 3.69e-19
C77 a_1108_47# a_1270_413# 0.006453f
C78 a_1108_47# a_543_47# 7.99e-20
C79 a_1217_47# a_1108_47# 0.007416f
C80 a_448_47# a_543_47# 0.049827f
C81 VGND RESET_B 0.287765f
C82 a_805_47# VGND 0.00579f
C83 a_639_47# a_543_47# 0.013793f
C84 VPB VPWR 0.21644f
C85 a_639_47# a_448_47# 4.61e-19
C86 a_1283_21# RESET_B 0.278137f
C87 a_651_413# a_761_289# 0.097745f
C88 VPWR D 0.081188f
C89 VPWR a_27_47# 0.152296f
C90 a_193_47# VPWR 0.395821f
C91 a_1108_47# RESET_B 0.236601f
C92 a_1270_413# RESET_B 2.06e-19
C93 VPB a_27_47# 0.261876f
C94 VPB D 0.137565f
C95 a_543_47# RESET_B 0.153272f
C96 a_448_47# RESET_B 2.45e-19
C97 VPB a_193_47# 0.17092f
C98 a_805_47# a_543_47# 0.001705f
C99 a_27_47# D 0.132849f
C100 a_1217_47# RESET_B 6.03e-19
C101 a_193_47# a_27_47# 0.906454f
C102 a_193_47# D 0.217945f
C103 a_639_47# RESET_B 9.54e-19
C104 Q VNB 0.089869f
C105 VGND VNB 1.02171f
C106 VPWR VNB 0.830843f
C107 RESET_B VNB 0.263863f
C108 D VNB 0.159894f
C109 CLK VNB 0.195254f
C110 VPB VNB 1.84511f
C111 a_651_413# VNB 0.004694f
C112 a_448_47# VNB 0.013901f
C113 a_1108_47# VNB 0.138544f
C114 a_1283_21# VNB 0.29898f
C115 a_543_47# VNB 0.157869f
C116 a_761_289# VNB 0.120848f
C117 a_193_47# VNB 0.273565f
C118 a_27_47# VNB 0.495775f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB a_75_212#
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
C0 X VGND 0.054484f
C1 a_75_212# VGND 0.104971f
C2 VGND VPB 0.005071f
C3 X VPWR 0.089604f
C4 a_75_212# VPWR 0.134042f
C5 VPWR VPB 0.035518f
C6 X A 8.48e-19
C7 a_75_212# A 0.177899f
C8 A VPB 0.052491f
C9 VPWR VGND 0.028869f
C10 VGND A 0.018424f
C11 VPWR A 0.021742f
C12 a_75_212# X 0.106512f
C13 X VPB 0.012788f
C14 a_75_212# VPB 0.057101f
C15 VGND VNB 0.20733f
C16 VPWR VNB 0.175531f
C17 X VNB 0.094159f
C18 A VNB 0.164205f
C19 VPB VNB 0.338976f
C20 a_75_212# VNB 0.210264f
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VPB VNB a_27_413# a_297_47# a_207_413#
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
C0 VGND X 0.065151f
C1 a_207_413# VPB 0.047771f
C2 VPWR A_N 0.018219f
C3 VPB B 0.111061f
C4 a_27_413# a_207_413# 0.185422f
C5 a_27_413# B 0.092611f
C6 a_207_413# a_297_47# 0.004764f
C7 VPWR X 0.055194f
C8 VPB A_N 0.080056f
C9 a_27_413# A_N 0.198147f
C10 X VPB 0.012221f
C11 a_207_413# B 0.181991f
C12 X a_297_47# 8.17e-20
C13 VGND VPWR 0.056424f
C14 a_207_413# A_N 8.2e-19
C15 VGND VPB 0.007626f
C16 VGND a_27_413# 0.086256f
C17 X a_207_413# 0.071579f
C18 VGND a_297_47# 0.005035f
C19 X B 0.030307f
C20 VPWR VPB 0.063352f
C21 VPWR a_27_413# 0.107953f
C22 VPWR a_297_47# 6.35e-19
C23 VGND a_207_413# 0.114823f
C24 VGND B 0.01869f
C25 a_27_413# VPB 0.083441f
C26 VPWR a_207_413# 0.111277f
C27 VGND A_N 0.047311f
C28 VPWR B 0.086692f
C29 VGND VNB 0.368472f
C30 X VNB 0.089221f
C31 VPWR VNB 0.291542f
C32 B VNB 0.132317f
C33 A_N VNB 0.201458f
C34 VPB VNB 0.604764f
C35 a_207_413# VNB 0.137402f
C36 a_27_413# VNB 0.196502f
.ends

.subckt sky130_fd_sc_hd__a31o_1 VPB VNB X A3 A2 A1 B1 VGND VPWR a_80_21# a_209_297#
+ a_209_47# a_303_47#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
C0 B1 VGND 0.017205f
C1 a_209_297# A2 0.036649f
C2 a_209_297# a_209_47# 6.96e-20
C3 a_209_297# a_80_21# 0.062574f
C4 VPB a_209_297# 0.002836f
C5 a_303_47# a_209_297# 1.26e-19
C6 A3 VGND 0.016898f
C7 A1 X 1.56e-19
C8 VPWR A1 0.018013f
C9 B1 a_80_21# 0.110759f
C10 VPB B1 0.034195f
C11 VGND X 0.057244f
C12 VPWR VGND 0.06622f
C13 A2 A3 0.108535f
C14 A3 a_209_47# 3.56e-19
C15 a_80_21# A3 0.116583f
C16 VPB A3 0.02968f
C17 A2 X 3.42e-19
C18 a_209_47# X 9.76e-19
C19 A2 VPWR 0.022678f
C20 VPWR a_209_47# 0.001019f
C21 a_80_21# X 0.076532f
C22 VPB X 0.010822f
C23 a_80_21# VPWR 0.09916f
C24 a_209_297# B1 0.006215f
C25 VPB VPWR 0.071542f
C26 a_303_47# X 6.01e-19
C27 a_303_47# VPWR 0.001051f
C28 VGND A1 0.013522f
C29 a_209_297# A3 0.02681f
C30 A2 A1 0.104261f
C31 a_80_21# A1 0.036671f
C32 a_209_297# VPWR 0.204727f
C33 VPB A1 0.028686f
C34 A2 VGND 0.014804f
C35 VGND a_209_47# 0.006958f
C36 a_80_21# VGND 0.216165f
C37 VPB VGND 0.007686f
C38 a_303_47# VGND 0.006612f
C39 B1 VPWR 0.01773f
C40 A2 a_80_21# 0.035741f
C41 A3 X 0.00625f
C42 a_209_297# A1 0.037771f
C43 a_80_21# a_209_47# 0.010132f
C44 VPB A2 0.028537f
C45 VPWR A3 0.040256f
C46 a_303_47# A2 3.38e-19
C47 VPB a_80_21# 0.050979f
C48 a_303_47# a_80_21# 0.011458f
C49 a_209_297# VGND 0.004304f
C50 VPWR X 0.117035f
C51 B1 A1 0.101116f
C52 VGND VNB 0.410332f
C53 VPWR VNB 0.331823f
C54 X VNB 0.08952f
C55 B1 VNB 0.11534f
C56 A1 VNB 0.089669f
C57 A2 VNB 0.089585f
C58 A3 VNB 0.089866f
C59 VPB VNB 0.69336f
C60 a_209_297# VNB 0.006211f
C61 a_80_21# VNB 0.211154f
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
C0 VPB VGND 0.161065f
C1 VPB VPWR 0.085759f
C2 VPWR VGND 0.903312f
C3 VPWR VNB 0.867393f
C4 VGND VNB 0.761362f
C5 VPB VNB 0.604764f
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 X A VPB VNB VGND VPWR a_49_47# a_285_47# a_391_47#
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
C0 a_285_47# VPB 0.156427f
C1 a_285_47# X 0.007197f
C2 a_285_47# VPWR 0.119832f
C3 a_49_47# a_391_47# 0.001885f
C4 a_285_47# A 0.001072f
C5 VGND a_285_47# 0.120945f
C6 VPB a_391_47# 0.044127f
C7 X a_391_47# 0.128943f
C8 VPWR a_391_47# 0.134775f
C9 VGND a_391_47# 0.130239f
C10 VPB a_49_47# 0.125413f
C11 VPWR a_49_47# 0.144268f
C12 VPB X 0.015496f
C13 a_49_47# A 0.279977f
C14 VGND a_49_47# 0.143546f
C15 VPWR VPB 0.0787f
C16 VPB A 0.082837f
C17 VGND VPB 0.007167f
C18 VPWR X 0.080229f
C19 a_285_47# a_391_47# 0.419086f
C20 VGND X 0.07961f
C21 VPWR A 0.020643f
C22 VGND VPWR 0.071507f
C23 VGND A 0.021393f
C24 a_285_47# a_49_47# 0.22264f
C25 VGND VNB 0.43965f
C26 X VNB 0.095447f
C27 VPWR VNB 0.367348f
C28 A VNB 0.178652f
C29 VPB VNB 0.781956f
C30 a_391_47# VNB 0.127705f
C31 a_285_47# VNB 0.29867f
C32 a_49_47# VNB 0.306903f
.ends

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VPB VNB a_561_47# a_297_297#
+ a_465_47# a_381_47# a_79_21#
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
C0 a_561_47# a_297_297# 3.62e-19
C1 X VPWR 0.063082f
C2 a_79_21# X 0.135998f
C3 VGND X 0.064052f
C4 X B1 1.21e-19
C5 a_297_297# A3 0.045547f
C6 a_297_297# A2 0.035373f
C7 a_381_47# a_297_297# 9.85e-19
C8 VPB A3 0.03038f
C9 a_297_297# VPWR 0.253629f
C10 a_297_297# A1 0.044438f
C11 A4 a_297_297# 0.03643f
C12 a_465_47# A3 0.001843f
C13 a_79_21# a_297_297# 0.053228f
C14 A2 VPB 0.027392f
C15 VGND a_297_297# 0.011109f
C16 a_465_47# A2 0.010642f
C17 VPB VPWR 0.081935f
C18 VPB A1 0.028093f
C19 A4 VPB 0.041818f
C20 a_79_21# VPB 0.052826f
C21 a_465_47# VPWR 8.18e-19
C22 VGND VPB 0.007308f
C23 B1 a_297_297# 0.002858f
C24 a_79_21# a_465_47# 5.59e-19
C25 VGND a_465_47# 0.004142f
C26 B1 VPB 0.043039f
C27 a_561_47# A3 0.009694f
C28 a_561_47# A2 9.72e-19
C29 X VPB 0.010526f
C30 a_561_47# VPWR 7.52e-19
C31 a_79_21# a_561_47# 2.93e-19
C32 VGND a_561_47# 0.006406f
C33 A2 A3 0.109547f
C34 a_381_47# A3 9.06e-20
C35 VPWR A3 0.024002f
C36 A3 A1 0.008128f
C37 A4 A3 0.108209f
C38 a_79_21# A3 6.62e-19
C39 a_297_297# VPB 0.006875f
C40 a_381_47# A2 0.008869f
C41 A2 VPWR 0.018762f
C42 VGND A3 0.074439f
C43 A2 A1 0.099595f
C44 a_465_47# a_297_297# 8.13e-19
C45 a_79_21# A2 0.030227f
C46 a_381_47# VPWR 8.83e-19
C47 a_381_47# A1 8.2e-20
C48 VGND A2 0.081373f
C49 VPWR A1 0.019035f
C50 A4 VPWR 0.020016f
C51 a_79_21# a_381_47# 0.002468f
C52 a_79_21# VPWR 0.124637f
C53 a_79_21# A1 0.008504f
C54 VGND a_381_47# 0.003407f
C55 a_79_21# A4 1.29e-19
C56 B1 A3 1.05e-19
C57 VGND VPWR 0.074653f
C58 VGND A1 0.016977f
C59 VGND A4 0.047952f
C60 a_79_21# VGND 0.144626f
C61 B1 A2 1.92e-19
C62 B1 VPWR 0.017677f
C63 B1 A1 0.099069f
C64 B1 A4 6.93e-21
C65 a_79_21# B1 0.149225f
C66 VGND B1 0.014254f
C67 VGND VNB 0.463871f
C68 VPWR VNB 0.364103f
C69 X VNB 0.092055f
C70 A4 VNB 0.156489f
C71 A3 VNB 0.099237f
C72 A2 VNB 0.096716f
C73 A1 VNB 0.093164f
C74 B1 VNB 0.112609f
C75 VPB VNB 0.781956f
C76 a_297_297# VNB 0.036501f
C77 a_79_21# VNB 0.141534f
.ends

.subckt sky130_fd_sc_hd__nor2_1 VPB VNB VGND VPWR A B Y a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 A Y 0.047068f
C1 A B 0.058413f
C2 VPWR A 0.052823f
C3 VGND VPB 0.004563f
C4 VGND Y 0.154448f
C5 VGND a_109_297# 0.001278f
C6 B VGND 0.045088f
C7 VPWR VGND 0.031443f
C8 Y VPB 0.013918f
C9 B VPB 0.036697f
C10 VPWR VPB 0.044857f
C11 Y a_109_297# 0.01129f
C12 B Y 0.087653f
C13 VPWR Y 0.099513f
C14 VPWR a_109_297# 0.006385f
C15 VPWR B 0.014836f
C16 A VGND 0.048556f
C17 A VPB 0.041461f
C18 VGND VNB 0.263197f
C19 VPWR VNB 0.214143f
C20 Y VNB 0.060508f
C21 A VNB 0.14927f
C22 B VNB 0.143121f
C23 VPB VNB 0.338976f
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
R1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
C0 VGND HI 0.206798f
C1 LO VGND 0.060475f
C2 VPB HI 0.004729f
C3 LO VPB 0.133883f
C4 VGND VPB 0.004789f
C5 VPWR HI 0.072643f
C6 VPWR LO 0.240897f
C7 VPWR VGND 0.031746f
C8 LO HI 0.068275f
C9 VPWR VPB 0.157853f
C10 VGND VNB 0.405957f
C11 LO VNB 0.165803f
C12 HI VNB 0.249567f
C13 VPWR VNB 0.297091f
C14 VPB VNB 0.338976f
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y a_199_47# a_113_297#
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
C0 Y A1 0.081255f
C1 Y a_113_297# 0.09093f
C2 VPB Y 0.014642f
C3 a_199_47# Y 0.001508f
C4 A1 B1 0.051837f
C5 B1 a_113_297# 0.007575f
C6 VPB B1 0.038865f
C7 A1 A2 0.091231f
C8 A2 a_113_297# 0.047625f
C9 A1 VPWR 0.015389f
C10 a_113_297# VPWR 0.1773f
C11 A1 VGND 0.077964f
C12 VPB A2 0.037282f
C13 VGND a_113_297# 0.008823f
C14 VPB VPWR 0.042396f
C15 VPB VGND 0.005478f
C16 a_199_47# VPWR 4.76e-19
C17 a_199_47# VGND 0.004279f
C18 Y B1 0.112603f
C19 Y A2 0.001218f
C20 Y VPWR 0.044654f
C21 Y VGND 0.065351f
C22 A1 a_113_297# 0.050014f
C23 B1 VPWR 0.01343f
C24 VPB A1 0.026387f
C25 VGND B1 0.043596f
C26 VPB a_113_297# 0.010797f
C27 a_199_47# A1 0.009167f
C28 a_199_47# a_113_297# 2.42e-19
C29 A2 VPWR 0.014703f
C30 A2 VGND 0.049477f
C31 VGND VPWR 0.036961f
C32 VGND VNB 0.285624f
C33 VPWR VNB 0.210674f
C34 Y VNB 0.054434f
C35 A2 VNB 0.143834f
C36 A1 VNB 0.098086f
C37 B1 VNB 0.161998f
C38 VPB VNB 0.427572f
C39 a_113_297# VNB 0.034004f
.ends

.subckt sky130_fd_sc_hd__o21a_1 VPB VNB VGND VPWR A1 A2 B1 X a_382_297# a_297_47#
+ a_79_21#
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VGND VPB 0.004903f
C1 VGND X 0.073624f
C2 VGND A2 0.017086f
C3 VPWR a_297_47# 0.005603f
C4 A1 VPB 0.041226f
C5 a_297_47# a_79_21# 0.032587f
C6 a_382_297# a_297_47# 8.13e-19
C7 A1 A2 0.102437f
C8 VPWR B1 0.021269f
C9 B1 a_79_21# 0.13448f
C10 VPWR VPB 0.062388f
C11 VPB a_79_21# 0.048932f
C12 X VPWR 0.095752f
C13 X a_79_21# 0.103737f
C14 A2 VPWR 0.083453f
C15 A2 a_79_21# 0.088854f
C16 VGND A1 0.015749f
C17 A2 a_382_297# 0.014523f
C18 a_297_47# B1 0.006369f
C19 a_297_47# VPB 7.6e-19
C20 VGND VPWR 0.058833f
C21 A2 a_297_47# 0.048027f
C22 VGND a_79_21# 0.129186f
C23 VGND a_382_297# 8.23e-19
C24 VPB B1 0.032789f
C25 X B1 3.56e-19
C26 A1 VPWR 0.044921f
C27 A1 a_79_21# 7.71e-19
C28 A2 B1 0.06645f
C29 A1 a_382_297# 2.25e-19
C30 X VPB 0.011001f
C31 A2 VPB 0.033371f
C32 VGND a_297_47# 0.124631f
C33 VPWR a_79_21# 0.201029f
C34 VPWR a_382_297# 0.00566f
C35 A1 a_297_47# 0.049229f
C36 a_382_297# a_79_21# 0.001446f
C37 VGND B1 0.018231f
C38 VGND VNB 0.351611f
C39 VPWR VNB 0.304004f
C40 X VNB 0.09354f
C41 A1 VNB 0.152087f
C42 A2 VNB 0.098105f
C43 B1 VNB 0.101193f
C44 VPB VNB 0.604764f
C45 a_297_47# VNB 0.034813f
C46 a_79_21# VNB 0.158207f
.ends

.subckt sky130_fd_sc_hd__inv_2 VPB VNB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 A VGND 0.063754f
C1 VGND Y 0.154601f
C2 VGND VPB 0.006491f
C3 VGND VPWR 0.042274f
C4 A Y 0.089386f
C5 A VPB 0.074183f
C6 A VPWR 0.06305f
C7 VPB Y 0.006097f
C8 Y VPWR 0.209105f
C9 VPB VPWR 0.052063f
C10 VGND VNB 0.266187f
C11 Y VNB 0.03316f
C12 VPWR VNB 0.246044f
C13 A VNB 0.262807f
C14 VPB VNB 0.338976f
.ends

.subckt r2r_dac_control VGND VPWR clk count[0] count[1] count[2] count[3] n_rst
XFILLER_0_13_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Left_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_27_ VGND VPWR VGND VPWR count[3] _04_ clknet_1_1__leaf_clk _27_/a_1020_47# _27_/a_975_413#
+ _27_/a_891_413# _27_/a_193_47# _27_/a_381_47# _27_/a_1062_300# _27_/a_572_47# _27_/a_568_413#
+ _27_/a_475_413# _27_/a_634_183# _27_/a_27_47# sky130_fd_sc_hd__dfxtp_4
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_55 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_26_ VGND VPWR VGND VPWR count[2] _03_ clknet_1_1__leaf_clk _26_/a_1020_47# _26_/a_975_413#
+ _26_/a_891_413# _26_/a_193_47# _26_/a_381_47# _26_/a_1062_300# _26_/a_572_47# _26_/a_568_413#
+ _26_/a_475_413# _26_/a_634_183# _26_/a_27_47# sky130_fd_sc_hd__dfxtp_4
XPHY_EDGE_ROW_1_Right_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25_ VGND VPWR VGND VPWR count[1] _02_ clknet_1_0__leaf_clk _25_/a_1020_47# _25_/a_975_413#
+ _25_/a_891_413# _25_/a_193_47# _25_/a_381_47# _25_/a_1062_300# _25_/a_572_47# _25_/a_568_413#
+ _25_/a_475_413# _25_/a_634_183# _25_/a_27_47# sky130_fd_sc_hd__dfxtp_4
XPHY_EDGE_ROW_7_Left_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk VGND VPWR VGND VPWR clk clknet_0_clk clkbuf_0_clk/a_110_47# sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24_ VGND VPWR VGND VPWR count[0] net4 clknet_1_0__leaf_clk _24_/a_1020_47# _24_/a_975_413#
+ _24_/a_891_413# _24_/a_193_47# _24_/a_381_47# _24_/a_1062_300# _24_/a_572_47# _24_/a_568_413#
+ _24_/a_475_413# _24_/a_634_183# _24_/a_27_47# sky130_fd_sc_hd__dfxtp_4
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23_ VGND VPWR VPWR VGND clknet_1_0__leaf_clk net2 _00_ rst _23_/a_1462_47# _23_/a_543_47#
+ _23_/a_651_413# _23_/a_193_47# _23_/a_805_47# _23_/a_448_47# _23_/a_639_47# _23_/a_1283_21#
+ _23_/a_761_289# _23_/a_1108_47# _23_/a_1217_47# _23_/a_1270_413# _23_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22_ VGND VPWR _04_ _10_ VPWR VGND _22_/a_75_212# sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21_ _10_ _08_ _09_ VGND VPWR VPWR VGND _21_/a_27_413# _21_/a_297_47# _21_/a_207_413#
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20_ VPWR VGND _09_ count[2] count[1] count[0] count[3] VGND VPWR _20_/a_80_21# _20_/a_209_297#
+ _20_/a_209_47# _20_/a_303_47# sky130_fd_sc_hd__a31o_1
Xinput1 VGND VPWR net1 n_rst VPWR VGND input1/a_75_212# sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_9_Right_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Right_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_89 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47#
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Right_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1 net3 rst VPWR VGND VGND VPWR hold1/a_49_47# hold1/a_285_47# hold1/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 net4 _01_ VPWR VGND VGND VPWR hold2/a_49_47# hold2/a_285_47# hold2/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19_ VGND VPWR count[2] count[3] count[1] _08_ rst count[0] VPWR VGND _19_/a_561_47#
+ _19_/a_297_297# _19_/a_465_47# _19_/a_381_47# _19_/a_79_21# sky130_fd_sc_hd__a41o_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 net5 count[2] VPWR VGND VGND VPWR hold3/a_49_47# hold3/a_285_47# hold3/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Left_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18_ VPWR VGND VGND VPWR _06_ _07_ _03_ _18_/a_109_297# sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_5_Left_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold4 net6 count[1] VPWR VGND VGND VPWR hold4/a_49_47# hold4/a_285_47# hold4/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17_ VPWR VGND _07_ count[2] count[1] count[0] net3 VGND VPWR _17_/a_80_21# _17_/a_209_297#
+ _17_/a_209_47# _17_/a_303_47# sky130_fd_sc_hd__a31o_1
XFILLER_0_15_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_15_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23__2 _23__2/LO net2 VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_16_ VPWR VGND VPWR VGND count[1] count[0] net5 _06_ _16_/a_199_47# _16_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47#
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15_ VPWR VGND VGND VPWR count[0] net6 _05_ _02_ _15_/a_382_297# _15_/a_297_47# _15_/a_79_21#
+ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_9_Left_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14_ VPWR VGND VPWR VGND count[1] count[0] net3 _05_ _14_/a_199_47# _14_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13_ VPWR VGND VGND VPWR count[0] net3 _01_ _13_/a_109_297# sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_7_Right_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12_ VPWR VGND VPWR VGND _00_ net1 sky130_fd_sc_hd__inv_2
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_13_Left_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_49 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Left_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
C0 _24_/a_193_47# net4 0.023423f
C1 _19_/a_297_297# _26_/a_27_47# 1.97e-19
C2 clknet_1_1__leaf_clk hold3/a_391_47# 3.86e-19
C3 net6 _25_/a_634_183# 2.13e-20
C4 net6 _24_/a_193_47# 0.383641f
C5 _22_/a_75_212# _27_/a_891_413# 6.62e-19
C6 _27_/a_572_47# clknet_0_clk 6.77e-19
C7 _20_/a_209_297# clkbuf_1_1__f_clk/a_110_47# 8.3e-20
C8 _23_/a_193_47# clk 9.45e-19
C9 hold1/a_391_47# _14_/a_113_297# 3.71e-19
C10 hold1/a_285_47# count[0] 0.02029f
C11 clknet_1_1__leaf_clk _06_ 0.001631f
C12 _23__2/LO _23_/a_27_47# 8.84e-20
C13 net6 _15_/a_382_297# 5.49e-19
C14 clknet_1_0__leaf_clk _23_/a_1283_21# 2.77e-19
C15 _21_/a_207_413# count[1] 7.99e-19
C16 clknet_1_0__leaf_clk count[2] 1.84e-20
C17 _21_/a_207_413# _27_/a_193_47# 2.32e-19
C18 _25_/a_572_47# count[1] 6.3e-20
C19 hold4/a_49_47# count[1] 0.064793f
C20 _25_/a_381_47# VPWR 0.002282f
C21 _26_/a_27_47# _20_/a_80_21# 2.47e-19
C22 net5 count[0] 0.005136f
C23 count[3] _27_/a_568_413# 0.001794f
C24 _26_/a_1062_300# count[0] 0.001057f
C25 _18_/a_109_297# count[0] 1.46e-19
C26 _08_ _22_/a_75_212# 2.09e-20
C27 clknet_1_0__leaf_clk _23_/a_543_47# 0.001108f
C28 _24_/a_475_413# VPWR -1.82e-19
C29 _01_ hold1/a_49_47# 8.61e-20
C30 _25_/a_975_413# clknet_1_0__leaf_clk 7.78e-19
C31 _20_/a_209_297# count[0] 0.002412f
C32 hold1/a_49_47# _24_/a_891_413# 7.62e-19
C33 _16_/a_113_297# VPWR 0.012564f
C34 _23__2/LO _15_/a_79_21# 4.17e-21
C35 _01_ count[1] 0.043335f
C36 _09_ _20_/a_209_297# 0.001922f
C37 clknet_1_0__leaf_clk _24_/a_1020_47# 4.93e-19
C38 hold1/a_49_47# VPWR 0.034542f
C39 _27_/a_27_47# clk 0.001076f
C40 _05_ _03_ 1.63e-20
C41 _07_ hold3/a_391_47# 0.027552f
C42 count[1] _24_/a_891_413# 0.002291f
C43 _26_/a_891_413# count[1] 0.001289f
C44 _24_/a_193_47# _24_/a_381_47# -0.008861f
C45 net3 _24_/a_475_413# 9.38e-21
C46 _03_ _17_/a_80_21# 5.14e-20
C47 count[1] VPWR 1.915105f
C48 _27_/a_193_47# VPWR 0.021204f
C49 hold2/a_285_47# rst 1.81e-19
C50 _23_/a_27_47# _24_/a_1062_300# 5.36e-20
C51 _23_/a_1108_47# _24_/a_1062_300# 0.002498f
C52 _27_/a_891_413# clk 3.4e-21
C53 count[3] _26_/a_975_413# 7.92e-20
C54 _25_/a_475_413# rst 2.67e-20
C55 count[3] rst 9.04e-19
C56 net3 _16_/a_113_297# 1.41e-19
C57 _07_ _06_ 0.017984f
C58 hold4/a_285_47# _24_/a_27_47# 6.76e-19
C59 net3 hold1/a_49_47# 0.020142f
C60 _17_/a_209_47# count[2] 0.00103f
C61 _16_/a_199_47# count[0] 0.001887f
C62 _25_/a_891_413# _24_/a_475_413# 0.001422f
C63 hold1/a_285_47# _25_/a_193_47# 1.77e-20
C64 _23_/a_761_289# clknet_0_clk 0.004317f
C65 net3 count[1] 0.250563f
C66 net1 _24_/a_891_413# 2.66e-21
C67 net2 VPWR 0.129689f
C68 _25_/a_1062_300# _01_ 1.71e-20
C69 _14_/a_113_297# count[2] 6.99e-20
C70 _08_ _06_ 8.98e-20
C71 clknet_1_1__leaf_clk net5 9.66e-19
C72 net1 VPWR 1.565992f
C73 _24_/a_193_47# clknet_0_clk 5.38e-20
C74 _25_/a_634_183# clknet_0_clk 1.53e-19
C75 clkbuf_0_clk/a_110_47# _24_/a_1062_300# 0.002632f
C76 hold1/a_391_47# _24_/a_475_413# 0.001791f
C77 clknet_1_1__leaf_clk _26_/a_1062_300# 6.12e-19
C78 _25_/a_1062_300# VPWR 0.032027f
C79 _15_/a_79_21# _24_/a_1062_300# 0.011454f
C80 _25_/a_891_413# count[1] 0.013219f
C81 clknet_1_1__leaf_clk _18_/a_109_297# 4.32e-19
C82 clknet_1_1__leaf_clk _20_/a_209_297# 0.001981f
C83 _19_/a_297_297# clknet_0_clk 0.001267f
C84 _00_ clk 4.3e-20
C85 _14_/a_199_47# count[1] 6.72e-19
C86 clknet_1_0__leaf_clk _24_/a_634_183# 0.037553f
C87 hold2/a_391_47# _24_/a_27_47# 5.09e-19
C88 _23_/a_1270_413# clknet_0_clk 2.2e-19
C89 _19_/a_465_47# count[1] 0.00215f
C90 _25_/a_475_413# clkbuf_1_0__f_clk/a_110_47# 0.007565f
C91 _21_/a_27_413# count[2] 0.001118f
C92 hold1/a_391_47# count[1] 0.025802f
C93 rst _04_ 2.78e-20
C94 hold3/a_49_47# count[0] 2.57e-19
C95 _23_/a_27_47# clkbuf_0_clk/a_110_47# 5.21e-20
C96 _25_/a_1062_300# net3 3.82e-19
C97 clknet_1_0__leaf_clk _23_/a_761_289# 7.87e-19
C98 _25_/a_1020_47# clknet_1_0__leaf_clk 6.14e-19
C99 _23__2/LO _23_/a_193_47# 8.84e-20
C100 clkbuf_0_clk/a_110_47# _19_/a_79_21# 0.00573f
C101 _20_/a_80_21# clknet_0_clk 0.00152f
C102 _25_/a_634_183# clknet_1_0__leaf_clk 0.034848f
C103 _15_/a_297_47# hold1/a_49_47# 0.038241f
C104 clknet_1_0__leaf_clk _24_/a_193_47# 0.432051f
C105 _26_/a_634_183# clkbuf_0_clk/a_110_47# 0.001372f
C106 _05_ _01_ 0.006259f
C107 _25_/a_27_47# _24_/a_891_413# 0.011052f
C108 _05_ _24_/a_891_413# 1.74e-21
C109 _07_ net5 0.107475f
C110 _25_/a_27_47# VPWR 0.069919f
C111 count[1] _15_/a_297_47# 2.36e-19
C112 count[0] _24_/a_1062_300# 0.068291f
C113 _03_ rst 9.87e-21
C114 _05_ VPWR 0.588812f
C115 count[3] _04_ 0.021904f
C116 _26_/a_891_413# _17_/a_80_21# 0.001212f
C117 _07_ _26_/a_1062_300# 0.0407f
C118 _25_/a_1062_300# hold1/a_391_47# 3.16e-20
C119 hold1/a_285_47# _24_/a_27_47# 5.81e-19
C120 hold4/a_391_47# count[1] 0.058649f
C121 _15_/a_79_21# clkbuf_0_clk/a_110_47# 0.008218f
C122 _17_/a_80_21# VPWR 0.079801f
C123 _17_/a_209_297# _24_/a_475_413# 1.16e-21
C124 _16_/a_113_297# _26_/a_193_47# 5.77e-20
C125 _08_ net5 4.85e-20
C126 hold4/a_285_47# net4 0.004768f
C127 hold1/a_49_47# _26_/a_193_47# 1.92e-21
C128 hold4/a_285_47# net6 0.002425f
C129 _26_/a_27_47# _06_ 4.35e-19
C130 hold3/a_285_47# count[3] 1.36e-20
C131 _25_/a_27_47# net3 2.79e-19
C132 _17_/a_209_297# hold1/a_49_47# 1.42e-20
C133 _24_/a_475_413# count[2] 1.46e-21
C134 _05_ net3 0.05478f
C135 count[1] _26_/a_193_47# 0.033958f
C136 _27_/a_193_47# _26_/a_193_47# 0.004458f
C137 _23_/a_27_47# count[0] 5.36e-20
C138 _23_/a_1108_47# count[0] 8.85e-19
C139 _17_/a_209_297# count[1] 5.06e-19
C140 net3 _17_/a_80_21# 0.016532f
C141 clknet_1_1__leaf_clk hold3/a_49_47# 2.47e-19
C142 _16_/a_113_297# count[2] 8.43e-19
C143 _08_ _20_/a_209_297# 5.19e-19
C144 _03_ count[3] 0.254623f
C145 _23_/a_193_47# _24_/a_1062_300# 2.17e-19
C146 _23_/a_1217_47# net2 7.68e-20
C147 hold2/a_391_47# _02_ 1.28e-19
C148 hold1/a_49_47# count[2] 5.75e-21
C149 _26_/a_475_413# clkbuf_0_clk/a_110_47# 0.001304f
C150 count[0] _19_/a_79_21# 0.012679f
C151 _26_/a_634_183# count[0] 0.019452f
C152 count[1] count[2] 0.244484f
C153 _07_ _16_/a_199_47# 3.04e-19
C154 _27_/a_193_47# count[2] 0.002804f
C155 _01_ _13_/a_109_297# 0.001105f
C156 _27_/a_568_413# VPWR -4.58e-19
C157 input1/a_75_212# _23_/a_27_47# 5.76e-20
C158 hold2/a_391_47# net4 0.002656f
C159 count[0] clkbuf_0_clk/a_110_47# 0.073435f
C160 net6 hold2/a_391_47# 1.2e-19
C161 _24_/a_193_47# _14_/a_113_297# 5.02e-20
C162 _09_ clkbuf_0_clk/a_110_47# 1.62e-21
C163 _15_/a_79_21# count[0] 0.002398f
C164 _13_/a_109_297# VPWR 6.8e-19
C165 _24_/a_975_413# VPWR 2.46e-19
C166 hold1/a_391_47# _17_/a_80_21# 5.26e-19
C167 _23_/a_27_47# _23_/a_193_47# -2.26e-19
C168 _17_/a_303_47# count[1] 0.00543f
C169 count[0] clkbuf_1_1__f_clk/a_110_47# 0.00143f
C170 net2 _23_/a_1283_21# 2.95e-20
C171 _25_/a_193_47# _24_/a_1062_300# 0.010477f
C172 net1 _23_/a_1283_21# 3.2e-19
C173 _25_/a_975_413# count[1] 6.67e-19
C174 _19_/a_561_47# count[0] 0.001203f
C175 hold1/a_285_47# _02_ 2.26e-19
C176 hold1/a_285_47# _26_/a_27_47# 2.16e-20
C177 _03_ _04_ 0.004737f
C178 count[1] _24_/a_1020_47# 2.72e-19
C179 _22_/a_75_212# clknet_0_clk 0.002695f
C180 _25_/a_27_47# _15_/a_297_47# 1.22e-20
C181 _01_ rst 0.001633f
C182 _21_/a_207_413# count[3] 2.1e-19
C183 _05_ _15_/a_297_47# 0.005004f
C184 net3 _24_/a_975_413# 5.13e-20
C185 net3 _13_/a_109_297# 0.001996f
C186 _07_ hold3/a_49_47# 0.001998f
C187 _23_/a_193_47# clkbuf_0_clk/a_110_47# 4.52e-20
C188 rst _24_/a_891_413# 1.27e-19
C189 _26_/a_475_413# count[0] 0.0249f
C190 net5 _26_/a_27_47# 0.001857f
C191 _23_/a_543_47# net2 0.002838f
C192 rst VPWR 0.760617f
C193 hold1/a_285_47# net4 0.002074f
C194 net1 _23_/a_543_47# 0.037397f
C195 net6 hold1/a_285_47# 1.83e-19
C196 hold3/a_285_47# _03_ 0.002726f
C197 _26_/a_572_47# count[0] 5.37e-19
C198 clknet_1_1__leaf_clk _19_/a_79_21# 2.84e-19
C199 _26_/a_1020_47# VPWR -4.44e-19
C200 _26_/a_634_183# clknet_1_1__leaf_clk 0.004487f
C201 _27_/a_475_413# clk 0.001919f
C202 _01_ hold2/a_285_47# 0.024954f
C203 _26_/a_27_47# _20_/a_209_297# 5.21e-20
C204 net3 rst 0.001416f
C205 clknet_1_1__leaf_clk clkbuf_0_clk/a_110_47# 0.001646f
C206 _26_/a_1062_300# net4 1.06e-21
C207 count[1] _26_/a_568_413# 2.02e-19
C208 _17_/a_80_21# _26_/a_193_47# 2.59e-20
C209 _25_/a_475_413# _24_/a_891_413# 0.001422f
C210 _26_/a_891_413# count[3] 4.33e-19
C211 hold2/a_285_47# VPWR 0.032704f
C212 _27_/a_27_47# _19_/a_79_21# 6.44e-19
C213 _25_/a_193_47# clkbuf_0_clk/a_110_47# 3.13e-20
C214 _25_/a_475_413# VPWR 0.006671f
C215 count[3] VPWR 2.360844f
C216 _10_ count[0] 8.84e-20
C217 _21_/a_27_413# _20_/a_80_21# 7.49e-20
C218 _21_/a_207_413# _04_ 3.53e-20
C219 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# 0.014091f
C220 _05_ count[2] 5.79e-19
C221 _10_ _09_ 0.002538f
C222 _24_/a_891_413# clkbuf_1_0__f_clk/a_110_47# 7.48e-19
C223 clknet_1_0__leaf_clk _24_/a_568_413# 4.58e-19
C224 _27_/a_27_47# clkbuf_0_clk/a_110_47# 7.77e-19
C225 _00_ _24_/a_1062_300# 9.63e-19
C226 VPWR clkbuf_1_0__f_clk/a_110_47# 0.111801f
C227 count[1] _24_/a_634_183# 0.007863f
C228 _17_/a_80_21# count[2] 0.041016f
C229 _24_/a_193_47# _24_/a_475_413# -0.021677f
C230 _23_/a_193_47# count[0] 1.16e-19
C231 net3 hold2/a_285_47# 0.001953f
C232 hold4/a_285_47# hold2/a_49_47# 0.001835f
C233 clk clknet_0_clk 0.037101f
C234 _19_/a_465_47# rst 4.82e-19
C235 n_rst VPWR 0.223836f
C236 net3 count[3] 1.66e-19
C237 hold1/a_391_47# rst 4.2e-19
C238 hold4/a_285_47# clknet_1_0__leaf_clk 0.006436f
C239 _25_/a_634_183# hold1/a_49_47# 2.83e-20
C240 hold1/a_49_47# _24_/a_193_47# 0.005676f
C241 clknet_1_1__leaf_clk _26_/a_475_413# 0.018417f
C242 _25_/a_1020_47# count[1] 7.25e-19
C243 _07_ _19_/a_79_21# 5.16e-20
C244 clknet_1_1__leaf_clk _26_/a_572_47# 0.001133f
C245 _23__2/LO _02_ 8.61e-20
C246 _26_/a_634_183# _07_ 0.001285f
C247 net3 clkbuf_1_0__f_clk/a_110_47# 2.02e-20
C248 _25_/a_634_183# count[1] 0.002382f
C249 _10_ _23_/a_193_47# 1.38e-20
C250 count[1] _24_/a_193_47# 0.057784f
C251 input1/a_75_212# _23_/a_193_47# 7.08e-20
C252 _00_ _23_/a_1108_47# 0.005452f
C253 _00_ _23_/a_27_47# 0.037394f
C254 count[0] _24_/a_572_47# 2.55e-19
C255 hold1/a_49_47# _15_/a_382_297# 2.23e-19
C256 _23_/a_1108_47# _24_/a_27_47# 3.63e-20
C257 clknet_1_1__leaf_clk count[0] 0.327982f
C258 _23_/a_27_47# _24_/a_27_47# 1.25e-19
C259 _04_ VPWR 0.304302f
C260 _08_ _19_/a_79_21# 0.005102f
C261 _25_/a_1062_300# _24_/a_634_183# 5.17e-19
C262 _15_/a_297_47# rst 0.004185f
C263 hold1/a_391_47# hold2/a_285_47# 3.65e-19
C264 clknet_1_1__leaf_clk _09_ 7.1e-19
C265 net2 _23_/a_761_289# 9.16e-19
C266 _25_/a_193_47# count[0] 0.030715f
C267 _25_/a_891_413# clkbuf_1_0__f_clk/a_110_47# 0.016063f
C268 _19_/a_297_297# count[1] 4.18e-19
C269 net1 _23_/a_761_289# 0.009364f
C270 _27_/a_381_47# clkbuf_0_clk/a_110_47# 4.3e-20
C271 _08_ clkbuf_0_clk/a_110_47# 0.00221f
C272 clknet_1_1__leaf_clk _10_ 6.95e-20
C273 clknet_1_0__leaf_clk hold2/a_391_47# 6.71e-19
C274 clknet_1_0__leaf_clk clk 1.7e-20
C275 hold3/a_285_47# VPWR 0.018853f
C276 _23_/a_1217_47# rst 1.58e-19
C277 _16_/a_113_297# _20_/a_80_21# 0.015784f
C278 _24_/a_27_47# clkbuf_0_clk/a_110_47# 2.46e-19
C279 _09_ _27_/a_27_47# 0.002125f
C280 _03_ _26_/a_891_413# 9.91e-20
C281 _25_/a_1062_300# _24_/a_193_47# 0.010477f
C282 _08_ clkbuf_1_1__f_clk/a_110_47# 3.08e-19
C283 _03_ VPWR 0.057985f
C284 count[1] _20_/a_80_21# 0.046236f
C285 _10_ _27_/a_27_47# 0.012996f
C286 count[3] _20_/a_209_47# 1.64e-20
C287 _07_ _26_/a_475_413# 1.54e-19
C288 _02_ _24_/a_1062_300# 0.024342f
C289 net1 _23_/a_1270_413# 1.04e-19
C290 _20_/a_209_297# clknet_0_clk 0.001397f
C291 _26_/a_975_413# count[2] 0.001258f
C292 _23_/a_1283_21# rst 0.019609f
C293 _25_/a_27_47# _24_/a_634_183# 8.67e-20
C294 _10_ _27_/a_891_413# 0.018642f
C295 _23_/a_805_47# clknet_0_clk 4.44e-19
C296 rst count[2] 0.009131f
C297 net3 _03_ 2.61e-20
C298 _07_ count[0] 0.03153f
C299 net4 _24_/a_1062_300# 3.52e-19
C300 clknet_1_0__leaf_clk hold1/a_285_47# 1.19e-19
C301 net6 _24_/a_1062_300# 0.053806f
C302 _23_/a_639_47# clknet_0_clk 7.29e-19
C303 _26_/a_1020_47# count[2] 7.75e-19
C304 count[3] _26_/a_193_47# 0.038233f
C305 _02_ _23_/a_1108_47# 0.001199f
C306 _02_ _23_/a_27_47# 5.51e-21
C307 _27_/a_1062_300# count[3] 0.065015f
C308 count[3] _17_/a_209_297# 6.38e-20
C309 _08_ count[0] 0.00186f
C310 _25_/a_27_47# _24_/a_193_47# 0.011266f
C311 _25_/a_27_47# _25_/a_634_183# -0.006998f
C312 _00_ count[0] 6.94e-19
C313 _23_/a_543_47# rst 2.05e-19
C314 _08_ _09_ 0.11537f
C315 _24_/a_27_47# count[0] 0.002154f
C316 clknet_1_1__leaf_clk _27_/a_27_47# 0.011461f
C317 _21_/a_297_47# VPWR -2.16e-19
C318 _21_/a_207_413# VPWR 0.011969f
C319 _25_/a_572_47# VPWR 2.52e-19
C320 hold4/a_49_47# VPWR 0.057951f
C321 _17_/a_80_21# _24_/a_193_47# 1.38e-20
C322 count[3] count[2] 0.504504f
C323 net6 _23_/a_1108_47# 2.38e-21
C324 net6 _23_/a_27_47# 5.8e-21
C325 _08_ _10_ 0.001045f
C326 _00_ _10_ 0.001743f
C327 _05_ _15_/a_382_297# 0.001001f
C328 _26_/a_27_47# clkbuf_0_clk/a_110_47# 9e-19
C329 clk _27_/a_634_183# 1.35e-19
C330 _02_ clkbuf_0_clk/a_110_47# 0.0039f
C331 clknet_1_1__leaf_clk _27_/a_891_413# 1.74e-19
C332 _23_/a_1217_47# _04_ 3.53e-21
C333 _23__2/LO clknet_0_clk 0.002049f
C334 _27_/a_975_413# count[3] 0.001926f
C335 _21_/a_27_413# _06_ 1.84e-20
C336 _15_/a_79_21# _02_ 0.034681f
C337 _26_/a_27_47# clkbuf_1_1__f_clk/a_110_47# 4.99e-19
C338 _00_ _23_/a_193_47# 0.03804f
C339 _26_/a_193_47# _04_ 1.85e-19
C340 _23_/a_193_47# _24_/a_27_47# 6.22e-21
C341 _27_/a_27_47# _27_/a_891_413# -0.001487f
C342 net6 clkbuf_0_clk/a_110_47# 0.010028f
C343 _01_ VPWR 0.563374f
C344 _19_/a_561_47# _02_ 1.61e-19
C345 clknet_1_1__leaf_clk _07_ 2.81e-19
C346 _27_/a_1062_300# _04_ 0.001508f
C347 _24_/a_891_413# VPWR -0.0018f
C348 _15_/a_79_21# net4 6.99e-20
C349 net6 _15_/a_79_21# 0.001639f
C350 _26_/a_891_413# VPWR 0.007841f
C351 _22_/a_75_212# count[1] 7.62e-20
C352 _22_/a_75_212# _27_/a_193_47# 0.001073f
C353 hold1/a_285_47# _14_/a_113_297# 0.002067f
C354 clknet_1_1__leaf_clk _27_/a_381_47# 2.4e-19
C355 _04_ count[2] 2.99e-19
C356 _26_/a_475_413# _26_/a_27_47# -0.001968f
C357 clknet_1_1__leaf_clk _08_ 0.00799f
C358 net3 _01_ 0.052629f
C359 count[1] _24_/a_568_413# 0.001097f
C360 net3 _24_/a_891_413# 3.84e-19
C361 net3 _26_/a_891_413# 7.7e-20
C362 _03_ _26_/a_193_47# 0.024095f
C363 _00_ _25_/a_193_47# 1.21e-19
C364 _24_/a_1062_300# clknet_0_clk 0.001325f
C365 net3 VPWR 0.447802f
C366 _26_/a_27_47# count[0] 0.05512f
C367 hold3/a_285_47# count[2] 0.027171f
C368 _25_/a_193_47# _24_/a_27_47# 0.011266f
C369 _02_ count[0] 0.126818f
C370 _27_/a_381_47# _27_/a_27_47# -0.008882f
C371 _08_ _27_/a_27_47# 0.037068f
C372 _26_/a_1062_300# _14_/a_113_297# 2.91e-21
C373 hold4/a_285_47# count[1] 0.069725f
C374 count[3] _26_/a_568_413# 3.97e-19
C375 rst _23_/a_761_289# 2.55e-19
C376 _16_/a_113_297# _06_ 0.009764f
C377 _03_ count[2] 0.017175f
C378 _25_/a_891_413# VPWR 0.002289f
C379 _27_/a_475_413# clkbuf_0_clk/a_110_47# 9.3e-20
C380 count[0] net4 0.002762f
C381 hold1/a_391_47# _01_ 2.42e-19
C382 net6 count[0] 0.197074f
C383 _25_/a_634_183# rst 3.5e-20
C384 rst _24_/a_193_47# 4.43e-20
C385 _26_/a_381_47# clkbuf_0_clk/a_110_47# 1.42e-19
C386 _14_/a_199_47# VPWR -4.35e-19
C387 count[1] _06_ 0.00909f
C388 _19_/a_465_47# VPWR -4.38e-19
C389 _23_/a_1108_47# clknet_0_clk 0.028697f
C390 _23_/a_27_47# clknet_0_clk 0.00939f
C391 hold1/a_391_47# VPWR -0.014904f
C392 _02_ _23_/a_193_47# 1.46e-20
C393 _15_/a_382_297# rst 0.002012f
C394 _25_/a_891_413# net3 3.86e-20
C395 _08_ _07_ 0.001481f
C396 _24_/a_634_183# clkbuf_1_0__f_clk/a_110_47# 8.64e-19
C397 clknet_0_clk _19_/a_79_21# 0.003388f
C398 count[1] hold2/a_391_47# 0.011259f
C399 clknet_1_0__leaf_clk _24_/a_1062_300# 0.010538f
C400 _26_/a_634_183# clknet_0_clk 2.25e-20
C401 _27_/a_193_47# clk 3.31e-20
C402 _07_ _24_/a_27_47# 5.88e-21
C403 net3 _14_/a_199_47# 0.001847f
C404 net3 hold1/a_391_47# 0.057411f
C405 clkbuf_0_clk/a_110_47# clknet_0_clk 0.173441f
C406 _08_ _27_/a_381_47# 0.008228f
C407 _15_/a_297_47# _24_/a_891_413# 6.63e-19
C408 _20_/a_209_47# VPWR 0.001711f
C409 _01_ hold4/a_391_47# 0.001525f
C410 _15_/a_297_47# VPWR -2.5e-19
C411 clknet_1_1__leaf_clk _02_ 9.54e-25
C412 clknet_1_1__leaf_clk _26_/a_27_47# 0.153501f
C413 hold1/a_285_47# _24_/a_475_413# 0.005182f
C414 _15_/a_79_21# clknet_0_clk 0.001079f
C415 _21_/a_297_47# count[2] 1.81e-19
C416 _21_/a_207_413# count[2] 0.001021f
C417 _24_/a_193_47# clkbuf_1_0__f_clk/a_110_47# 9.68e-19
C418 _25_/a_634_183# clkbuf_1_0__f_clk/a_110_47# 0.006568f
C419 net2 clk 3.74e-20
C420 _00_ _24_/a_27_47# 6.3e-20
C421 clknet_0_clk clkbuf_1_1__f_clk/a_110_47# 0.013268f
C422 _02_ _25_/a_193_47# 0.041984f
C423 hold4/a_391_47# VPWR 0.03375f
C424 _23_/a_651_413# _23_/a_193_47# -0.007045f
C425 _25_/a_891_413# hold1/a_391_47# 3.49e-19
C426 net1 clk 0.001113f
C427 _19_/a_297_297# count[3] 0.01079f
C428 _23_/a_1217_47# VPWR 1.22e-19
C429 clknet_1_0__leaf_clk _23_/a_1108_47# 1.14e-19
C430 clknet_1_0__leaf_clk _23_/a_27_47# 0.018772f
C431 count[0] _24_/a_381_47# 1.06e-19
C432 _09_ _27_/a_475_413# 2.8e-19
C433 net6 _24_/a_572_47# 0.001444f
C434 _26_/a_381_47# count[0] 2.64e-19
C435 _25_/a_1062_300# hold2/a_391_47# 0.001063f
C436 _27_/a_27_47# _26_/a_27_47# 0.076413f
C437 _26_/a_891_413# _26_/a_193_47# -0.001f
C438 hold1/a_285_47# count[1] 0.017587f
C439 _26_/a_193_47# VPWR 0.003918f
C440 net6 _25_/a_193_47# 8.6e-19
C441 _10_ _27_/a_475_413# 0.001281f
C442 _27_/a_1062_300# VPWR 0.065824f
C443 _26_/a_475_413# clknet_0_clk 4.58e-20
C444 _17_/a_209_297# VPWR 1.3e-19
C445 _01_ count[2] 0.001917f
C446 count[3] _20_/a_80_21# 0.016094f
C447 clknet_1_0__leaf_clk clkbuf_0_clk/a_110_47# 0.001048f
C448 net5 count[1] 8.94e-19
C449 _10_ _20_/a_303_47# 1.78e-19
C450 _26_/a_891_413# count[2] 0.049539f
C451 _16_/a_113_297# _20_/a_209_297# 4.94e-20
C452 _23_/a_1283_21# VPWR 0.044416f
C453 _26_/a_1062_300# count[1] 1.01e-19
C454 VPWR count[2] 1.623981f
C455 net3 _26_/a_193_47# 4.27e-19
C456 count[0] clknet_0_clk 0.179312f
C457 _05_ _06_ 2.1e-20
C458 net3 _17_/a_209_297# 5.3e-20
C459 _09_ clknet_0_clk 0.010726f
C460 _07_ _26_/a_27_47# 5.44e-19
C461 count[1] _20_/a_209_297# 0.03427f
C462 _27_/a_975_413# VPWR -2.85e-19
C463 _17_/a_80_21# _06_ 5.3e-21
C464 _17_/a_303_47# VPWR -0.001051f
C465 _10_ clknet_0_clk 0.139387f
C466 net3 count[2] 0.079424f
C467 _05_ clk 2.08e-19
C468 _27_/a_381_47# _26_/a_27_47# 4.83e-21
C469 _23_/a_543_47# VPWR 0.018102f
C470 clknet_1_1__leaf_clk _27_/a_475_413# 1.88e-19
C471 _08_ _26_/a_27_47# 0.005307f
C472 _00_ _02_ 0.001234f
C473 _27_/a_572_47# VPWR 2.67e-19
C474 _24_/a_1020_47# VPWR -2.83e-19
C475 clknet_1_1__leaf_clk _26_/a_381_47# 0.010653f
C476 _02_ _24_/a_27_47# 5.09e-20
C477 _23_/a_193_47# clknet_0_clk 0.012059f
C478 _03_ _15_/a_382_297# 6.5e-20
C479 net2 _23_/a_805_47# 4.48e-19
C480 hold2/a_49_47# count[0] 1.8e-19
C481 _17_/a_303_47# net3 9.02e-19
C482 _03_ _19_/a_297_297# 3.25e-19
C483 _27_/a_27_47# _27_/a_475_413# -0.026874f
C484 clknet_1_0__leaf_clk count[0] 0.50536f
C485 _22_/a_75_212# rst 2.96e-21
C486 _23_/a_639_47# net2 0.001136f
C487 _24_/a_27_47# net4 0.039287f
C488 hold3/a_285_47# _20_/a_80_21# 1.3e-19
C489 _23_/a_1462_47# clknet_0_clk 6.77e-19
C490 net6 _24_/a_27_47# 0.035053f
C491 _26_/a_381_47# _27_/a_27_47# 4.83e-21
C492 _25_/a_27_47# hold1/a_285_47# 8.16e-21
C493 _05_ hold1/a_285_47# 0.00102f
C494 _03_ _20_/a_80_21# 0.018221f
C495 clknet_1_1__leaf_clk clknet_0_clk 0.031819f
C496 _00_ _23_/a_651_413# 0.001582f
C497 input1/a_75_212# clknet_1_0__leaf_clk 0.001023f
C498 _25_/a_193_47# clknet_0_clk 0.001434f
C499 hold1/a_285_47# _17_/a_80_21# 2.56e-20
C500 _25_/a_381_47# _24_/a_1062_300# 5.68e-19
C501 hold4/a_49_47# _24_/a_193_47# 2.17e-19
C502 VPWR _26_/a_568_413# 1.67e-19
C503 _21_/a_27_413# _19_/a_79_21# 1.44e-21
C504 clknet_1_0__leaf_clk _23_/a_193_47# 0.007442f
C505 _20_/a_209_47# count[2] 0.004735f
C506 _22_/a_75_212# count[3] 9.86e-20
C507 _27_/a_27_47# clknet_0_clk 0.02579f
C508 _17_/a_80_21# net5 7.13e-22
C509 _27_/a_1020_47# _10_ 7.77e-19
C510 _21_/a_27_413# clkbuf_0_clk/a_110_47# 1.03e-19
C511 _24_/a_634_183# VPWR 0.004977f
C512 _26_/a_1062_300# _17_/a_80_21# 3.58e-19
C513 _27_/a_891_413# clknet_0_clk 6.1e-19
C514 _17_/a_209_297# _26_/a_193_47# 2.21e-19
C515 _08_ _27_/a_475_413# 0.005988f
C516 hold1/a_49_47# _24_/a_1062_300# 8.33e-19
C517 _23_/a_761_289# VPWR 0.022066f
C518 count[1] _24_/a_1062_300# 8.04e-19
C519 _24_/a_27_47# _24_/a_381_47# -0.005913f
C520 _08_ _20_/a_303_47# 7.49e-19
C521 _26_/a_193_47# count[2] 0.046072f
C522 _25_/a_634_183# _24_/a_891_413# 0.001115f
C523 hold2/a_391_47# rst 1.37e-19
C524 clknet_1_0__leaf_clk _25_/a_193_47# 0.229333f
C525 net3 _24_/a_634_183# 5.4e-21
C526 _25_/a_634_183# VPWR 0.00743f
C527 rst clk 0.005073f
C528 count[0] _14_/a_113_297# 0.045104f
C529 _24_/a_193_47# VPWR -0.001592f
C530 _17_/a_209_297# count[2] 0.033969f
C531 _19_/a_381_47# count[0] 0.00285f
C532 _01_ _15_/a_382_297# 1.03e-21
C533 _02_ net4 1.1e-19
C534 net6 _26_/a_27_47# 9.87e-21
C535 net6 _02_ 0.082646f
C536 _22_/a_75_212# _04_ 0.002083f
C537 count[3] _06_ 8.29e-20
C538 _15_/a_382_297# VPWR 2.64e-19
C539 _27_/a_381_47# clknet_0_clk 0.004027f
C540 _25_/a_891_413# _24_/a_634_183# 0.001115f
C541 _19_/a_297_297# VPWR 0.061473f
C542 _08_ clknet_0_clk 0.115145f
C543 _23_/a_193_47# _23_/a_448_47# -0.004818f
C544 net1 _24_/a_1062_300# 8.73e-20
C545 net3 _25_/a_634_183# 1.29e-19
C546 net3 _24_/a_193_47# 0.001882f
C547 _23_/a_1270_413# VPWR 7.02e-20
C548 net6 net4 0.028023f
C549 _00_ clknet_0_clk 0.135559f
C550 _10_ _27_/a_634_183# 0.009529f
C551 _26_/a_634_183# _16_/a_113_297# 6.18e-20
C552 _24_/a_27_47# clknet_0_clk 4.22e-20
C553 _23__2/LO _05_ 5.95e-22
C554 _26_/a_634_183# hold1/a_49_47# 8.55e-21
C555 hold1/a_391_47# _24_/a_634_183# 4.06e-19
C556 count[3] clk 0.15287f
C557 _17_/a_303_47# count[2] 1.8e-19
C558 _21_/a_27_413# _09_ 0.095071f
C559 count[1] _19_/a_79_21# 0.003341f
C560 _27_/a_193_47# _19_/a_79_21# 4.32e-19
C561 net3 _15_/a_382_297# 1.94e-19
C562 _26_/a_634_183# count[1] 0.002701f
C563 _25_/a_891_413# _24_/a_193_47# 5.66e-20
C564 hold1/a_285_47# rst 0.00209f
C565 hold1/a_49_47# clkbuf_0_clk/a_110_47# 0.01619f
C566 _20_/a_80_21# VPWR 0.03208f
C567 _21_/a_27_413# _10_ 4.68e-19
C568 _15_/a_79_21# hold1/a_49_47# 0.001296f
C569 count[1] clkbuf_0_clk/a_110_47# 0.007577f
C570 _23_/a_27_47# net2 0.041949f
C571 _23_/a_1108_47# net2 6.62e-19
C572 _27_/a_193_47# clkbuf_0_clk/a_110_47# 9.44e-20
C573 net1 _23_/a_1108_47# 0.002028f
C574 n_rst clk 0.050543f
C575 net1 _23_/a_27_47# 0.051346f
C576 hold1/a_391_47# _24_/a_193_47# 0.005482f
C577 count[1] clkbuf_1_1__f_clk/a_110_47# 0.001171f
C578 _25_/a_381_47# count[0] 0.004498f
C579 _26_/a_381_47# _26_/a_27_47# -0.005059f
C580 _00_ clknet_1_0__leaf_clk 0.06156f
C581 hold2/a_285_47# hold1/a_285_47# 0.005423f
C582 clknet_1_1__leaf_clk _27_/a_634_183# 1.82e-19
C583 _19_/a_561_47# count[1] 0.002728f
C584 clknet_1_0__leaf_clk _24_/a_27_47# 0.271496f
C585 _16_/a_113_297# _26_/a_475_413# 1.39e-19
C586 _03_ hold3/a_391_47# 8.59e-19
C587 _23_/a_805_47# rst 1.11e-19
C588 _25_/a_27_47# _24_/a_1062_300# 0.004485f
C589 _04_ clk 1.2e-19
C590 hold3/a_285_47# _06_ 0.001413f
C591 _05_ _24_/a_1062_300# 0.011659f
C592 net4 _24_/a_381_47# 0.007326f
C593 count[0] _24_/a_475_413# 0.001299f
C594 hold1/a_285_47# clkbuf_1_0__f_clk/a_110_47# 2e-21
C595 net6 _24_/a_381_47# 0.014464f
C596 _25_/a_568_413# VPWR 3.1e-19
C597 count[1] _26_/a_475_413# 0.012159f
C598 net6 _26_/a_381_47# 1.08e-19
C599 _27_/a_27_47# _27_/a_634_183# -0.012442f
C600 _23_/a_639_47# rst 1.76e-19
C601 _26_/a_568_413# count[2] 1.6e-19
C602 clknet_1_1__leaf_clk _21_/a_27_413# 3.86e-19
C603 _26_/a_572_47# count[1] 1.15e-19
C604 _03_ _06_ 0.043866f
C605 _16_/a_113_297# count[0] 0.047081f
C606 hold4/a_391_47# _24_/a_193_47# 7.18e-19
C607 count[3] _26_/a_1062_300# 2.99e-19
C608 hold1/a_49_47# count[0] 0.041094f
C609 _02_ clknet_0_clk 0.038218f
C610 _26_/a_27_47# clknet_0_clk 4.09e-20
C611 count[1] count[0] 1.640845f
C612 count[3] _20_/a_209_297# 2.24e-20
C613 _21_/a_27_413# _27_/a_27_47# 0.010277f
C614 _09_ count[1] 0.008704f
C615 _09_ _27_/a_193_47# 0.008413f
C616 _17_/a_209_297# _24_/a_193_47# 1.02e-20
C617 net6 clknet_0_clk 0.001818f
C618 _23__2/LO rst 7.45e-20
C619 _10_ count[1] 2.57e-19
C620 _00_ _23_/a_448_47# 5.52e-19
C621 _10_ _27_/a_193_47# 0.022613f
C622 _23_/a_1283_21# _24_/a_193_47# 6.57e-20
C623 _24_/a_193_47# count[2] 3.07e-21
C624 net1 count[0] 0.001688f
C625 _25_/a_27_47# clkbuf_0_clk/a_110_47# 4.23e-19
C626 _26_/a_634_183# _17_/a_80_21# 6.22e-20
C627 _25_/a_381_47# _25_/a_193_47# -0.001414f
C628 _05_ clkbuf_0_clk/a_110_47# 0.045833f
C629 hold2/a_49_47# _02_ 7.32e-21
C630 _22_/a_75_212# VPWR 0.068177f
C631 _08_ _27_/a_634_183# 0.001694f
C632 _21_/a_207_413# _06_ 3.21e-20
C633 _25_/a_27_47# _15_/a_79_21# 2.97e-19
C634 clknet_1_0__leaf_clk _02_ 0.082338f
C635 _24_/a_27_47# _14_/a_113_297# 6.97e-20
C636 _25_/a_1062_300# count[0] 2.79e-20
C637 _17_/a_80_21# clkbuf_0_clk/a_110_47# 0.001119f
C638 _15_/a_79_21# _05_ 0.031226f
C639 _24_/a_568_413# VPWR 2.87e-20
C640 hold3/a_285_47# net5 0.001274f
C641 _19_/a_297_297# count[2] 0.013553f
C642 input1/a_75_212# net2 3.23e-19
C643 hold4/a_285_47# _01_ 0.001434f
C644 clknet_1_1__leaf_clk _16_/a_113_297# 0.005869f
C645 hold2/a_49_47# net4 0.001341f
C646 input1/a_75_212# net1 0.001973f
C647 net6 hold2/a_49_47# 0.004417f
C648 clknet_1_0__leaf_clk net4 0.078761f
C649 _21_/a_27_413# _27_/a_381_47# 8.01e-19
C650 hold3/a_285_47# _26_/a_1062_300# 0.021006f
C651 net6 clknet_1_0__leaf_clk 0.132677f
C652 count[1] _24_/a_572_47# 5.42e-19
C653 hold4/a_285_47# VPWR 0.044492f
C654 _21_/a_27_413# _08_ 0.025245f
C655 _03_ net5 0.267742f
C656 _23_/a_193_47# net2 1.17e-19
C657 net1 _23_/a_193_47# 0.424952f
C658 clknet_1_1__leaf_clk count[1] 0.334917f
C659 hold3/a_285_47# _20_/a_209_297# 4.92e-20
C660 clknet_1_1__leaf_clk _27_/a_193_47# 0.001808f
C661 _27_/a_475_413# clknet_0_clk 0.015559f
C662 VPWR hold3/a_391_47# 0.007567f
C663 _03_ _26_/a_1062_300# 6e-19
C664 count[1] _25_/a_193_47# 0.004001f
C665 _20_/a_80_21# count[2] 0.05524f
C666 rst _24_/a_1062_300# 0.008392f
C667 clknet_1_0__leaf_clk _23_/a_651_413# 8.11e-19
C668 _26_/a_891_413# _06_ 5.84e-19
C669 _17_/a_80_21# _26_/a_475_413# 0.001305f
C670 VPWR _06_ 0.132711f
C671 _25_/a_27_47# count[0] 0.02934f
C672 _27_/a_193_47# _27_/a_27_47# -0.116315f
C673 _01_ hold2/a_391_47# 0.009007f
C674 _05_ count[0] 0.210006f
C675 _17_/a_80_21# count[0] 0.046062f
C676 net1 _25_/a_193_47# 9.22e-20
C677 clk VPWR 0.672313f
C678 hold2/a_391_47# VPWR 0.016085f
C679 _00_ _25_/a_381_47# 5.08e-20
C680 _23_/a_1108_47# rst 0.001344f
C681 _23_/a_27_47# rst 1.76e-19
C682 _25_/a_475_413# _24_/a_1062_300# 0.007354f
C683 net3 _06_ 2.63e-21
C684 _03_ _16_/a_199_47# 7.25e-19
C685 rst _19_/a_79_21# 0.050697f
C686 _24_/a_1062_300# clkbuf_1_0__f_clk/a_110_47# 0.002145f
C687 clknet_1_0__leaf_clk _24_/a_381_47# 0.013889f
C688 _07_ count[1] 0.055679f
C689 _24_/a_27_47# _24_/a_475_413# -0.006348f
C690 _24_/a_193_47# _24_/a_634_183# -0.013106f
C691 net3 clk 0.001347f
C692 net3 hold2/a_391_47# 0.006395f
C693 _08_ _16_/a_113_297# 1.69e-19
C694 rst clkbuf_0_clk/a_110_47# 0.067245f
C695 _01_ hold1/a_285_47# 2.96e-19
C696 _27_/a_381_47# _27_/a_193_47# -0.001414f
C697 hold1/a_49_47# _24_/a_27_47# 0.010568f
C698 _15_/a_79_21# rst 0.06472f
C699 _26_/a_891_413# hold1/a_285_47# 4.26e-20
C700 _08_ count[1] 0.002618f
C701 _08_ _27_/a_193_47# 0.042353f
C702 hold1/a_285_47# VPWR -0.0135f
C703 count[1] _24_/a_27_47# 0.277438f
C704 _25_/a_634_183# _24_/a_193_47# 8.84e-20
C705 count[3] _19_/a_79_21# 4.73e-19
C706 clknet_1_0__leaf_clk clknet_0_clk 0.045368f
C707 _19_/a_561_47# rst 3.85e-19
C708 _26_/a_634_183# count[3] 4.49e-19
C709 _27_/a_1062_300# _22_/a_75_212# 3.46e-19
C710 count[0] _24_/a_975_413# 3.96e-19
C711 _13_/a_109_297# count[0] 9.92e-21
C712 _26_/a_891_413# net5 5.4e-19
C713 _03_ hold3/a_49_47# 4.56e-19
C714 _25_/a_27_47# _25_/a_193_47# -0.135024f
C715 hold1/a_391_47# hold2/a_391_47# 0.009581f
C716 net5 VPWR 0.033453f
C717 n_rst _23_/a_27_47# 0.002092f
C718 _05_ _25_/a_193_47# 4.09e-20
C719 count[3] clkbuf_0_clk/a_110_47# 0.009679f
C720 _25_/a_475_413# clkbuf_0_clk/a_110_47# 4.17e-19
C721 net3 hold1/a_285_47# 0.081218f
C722 _00_ net2 0.010695f
C723 _22_/a_75_212# count[2] 5.65e-21
C724 _26_/a_1062_300# VPWR 0.014942f
C725 _00_ net1 0.132167f
C726 _18_/a_109_297# VPWR 1.28e-19
C727 count[3] clkbuf_1_1__f_clk/a_110_47# 4.25e-19
C728 _20_/a_209_297# VPWR 0.005733f
C729 _02_ _25_/a_381_47# 0.004581f
C730 _26_/a_975_413# count[0] 4.79e-19
C731 net3 net5 2.24e-21
C732 _23_/a_1108_47# _04_ 4.08e-20
C733 rst count[0] 0.299439f
C734 _25_/a_1062_300# _24_/a_27_47# 0.004485f
C735 _23_/a_27_47# _04_ 6.27e-23
C736 net3 _26_/a_1062_300# 3.31e-21
C737 _09_ rst 1.75e-20
C738 _23_/a_639_47# VPWR 8.89e-20
C739 _04_ _19_/a_79_21# 1.09e-20
C740 _26_/a_1020_47# count[0] 5.16e-19
C741 _26_/a_193_47# _06_ 3.98e-19
C742 count[3] _26_/a_475_413# 0.003068f
C743 hold3/a_391_47# count[2] 0.011804f
C744 _17_/a_209_297# _06_ 3.86e-20
C745 _10_ rst 0.003632f
C746 _16_/a_113_297# _26_/a_27_47# 8.02e-20
C747 hold1/a_49_47# _26_/a_27_47# 2.56e-21
C748 hold1/a_49_47# _02_ 0.001005f
C749 _04_ clkbuf_0_clk/a_110_47# 0.003431f
C750 _16_/a_199_47# VPWR -3.11e-19
C751 _23_/a_448_47# clknet_0_clk 4.34e-19
C752 hold2/a_285_47# count[0] 3.51e-19
C753 net4 _24_/a_475_413# 0.001175f
C754 _21_/a_27_413# _27_/a_475_413# 1.23e-20
C755 net6 _24_/a_475_413# 0.02387f
C756 count[1] _02_ 1.45e-19
C757 count[1] _26_/a_27_47# 0.030415f
C758 count[3] count[0] 0.070048f
C759 _07_ _17_/a_80_21# 0.001652f
C760 _06_ count[2] 0.003864f
C761 _25_/a_475_413# count[0] 0.017906f
C762 _27_/a_193_47# _26_/a_27_47# 7.18e-19
C763 _23_/a_193_47# rst 1.95e-19
C764 _09_ count[3] 6.81e-19
C765 hold1/a_391_47# _26_/a_1062_300# 3.58e-20
C766 hold1/a_49_47# net4 4.16e-19
C767 _27_/a_27_47# _27_/a_568_413# -9.71e-19
C768 _00_ _25_/a_27_47# 1.86e-19
C769 _23__2/LO VPWR 0.13462f
C770 net6 hold1/a_49_47# 0.006534f
C771 clknet_0_clk _27_/a_634_183# 0.01188f
C772 count[0] clkbuf_1_0__f_clk/a_110_47# 0.05437f
C773 _26_/a_634_183# _03_ 6.62e-19
C774 _25_/a_27_47# _24_/a_27_47# 0.001547f
C775 net3 _16_/a_199_47# 9.58e-20
C776 _23_/a_1283_21# clk 0.001675f
C777 _05_ _24_/a_27_47# 5.85e-21
C778 _08_ _17_/a_80_21# 8.13e-20
C779 count[1] net4 0.132658f
C780 _23_/a_1462_47# rst 8.75e-19
C781 net6 count[1] 0.079635f
C782 _10_ count[3] 0.035414f
C783 _03_ clkbuf_0_clk/a_110_47# 0.001063f
C784 _02_ net2 5.95e-22
C785 _17_/a_80_21# _24_/a_27_47# 1.15e-20
C786 net1 _02_ 0.001884f
C787 clknet_1_1__leaf_clk rst 0.00839f
C788 hold3/a_49_47# VPWR 0.066515f
C789 _21_/a_27_413# clknet_0_clk 0.005931f
C790 _03_ clkbuf_1_1__f_clk/a_110_47# 3.06e-19
C791 clknet_1_0__leaf_clk _23_/a_448_47# 0.001272f
C792 _25_/a_1062_300# _02_ 3.4e-19
C793 hold1/a_285_47# _17_/a_209_297# 2.44e-20
C794 n_rst input1/a_75_212# 0.02012f
C795 _04_ count[0] 4.42e-20
C796 _27_/a_27_47# rst 0.00168f
C797 _09_ _04_ 1.13e-20
C798 net5 _26_/a_193_47# 0.009094f
C799 n_rst _23_/a_193_47# 4.1e-19
C800 _25_/a_1062_300# net4 0.013058f
C801 _25_/a_1062_300# net6 6.02e-20
C802 hold1/a_285_47# count[2] 5.89e-19
C803 _03_ _26_/a_475_413# 0.002274f
C804 _24_/a_1062_300# VPWR 0.017331f
C805 _08_ _27_/a_568_413# 5.17e-19
C806 _26_/a_1062_300# _26_/a_193_47# -0.001214f
C807 hold3/a_285_47# count[0] 9.98e-19
C808 clknet_1_1__leaf_clk count[3] 0.067521f
C809 net1 _23_/a_651_413# 0.031249f
C810 _10_ _04_ 0.154238f
C811 _26_/a_1062_300# _17_/a_209_297# 5.78e-19
C812 hold3/a_285_47# _09_ 8.63e-21
C813 _25_/a_381_47# clknet_0_clk 2.89e-19
C814 _25_/a_475_413# _25_/a_193_47# -0.003996f
C815 net5 count[2] 0.003824f
C816 _27_/a_193_47# _27_/a_475_413# -0.003996f
C817 count[1] _24_/a_381_47# 0.021987f
C818 _03_ count[0] 0.185566f
C819 _26_/a_381_47# count[1] 0.004185f
C820 _26_/a_1062_300# count[2] 0.113922f
C821 _25_/a_193_47# clkbuf_1_0__f_clk/a_110_47# 0.011307f
C822 count[3] _27_/a_27_47# 0.42738f
C823 _25_/a_27_47# _02_ 0.017015f
C824 _07_ rst 2.41e-20
C825 _18_/a_109_297# count[2] 5.61e-19
C826 _05_ _02_ 0.11331f
C827 _05_ _26_/a_27_47# 6.62e-21
C828 _23_/a_27_47# _24_/a_891_413# 1.11e-20
C829 _23_/a_27_47# VPWR 0.039205f
C830 _23_/a_1108_47# VPWR 0.021961f
C831 _20_/a_209_297# count[2] 0.006947f
C832 hold4/a_285_47# _24_/a_193_47# 2.99e-19
C833 count[3] _27_/a_891_413# 0.039874f
C834 _17_/a_80_21# _26_/a_27_47# 6.11e-20
C835 _07_ _26_/a_1020_47# 7.13e-19
C836 hold1/a_49_47# clknet_0_clk 0.002956f
C837 net6 _25_/a_27_47# 2.74e-19
C838 VPWR _19_/a_79_21# 0.061565f
C839 _08_ rst 0.052447f
C840 _05_ net4 3.55e-20
C841 _01_ clkbuf_0_clk/a_110_47# 9.06e-20
C842 _00_ rst 4.99e-19
C843 net6 _05_ 0.076184f
C844 _26_/a_634_183# VPWR 0.008052f
C845 clknet_1_1__leaf_clk _04_ 0.002367f
C846 rst _24_/a_27_47# 6.23e-20
C847 count[1] clknet_0_clk 0.0109f
C848 clkbuf_0_clk/a_110_47# _24_/a_891_413# 8.66e-19
C849 _27_/a_193_47# clknet_0_clk 0.03508f
C850 _15_/a_79_21# _01_ 2.11e-21
C851 clknet_1_0__leaf_clk _25_/a_381_47# 0.013966f
C852 _25_/a_1062_300# _24_/a_381_47# 5.68e-19
C853 _07_ count[3] 9.8e-20
C854 clkbuf_0_clk/a_110_47# VPWR 0.169876f
C855 _15_/a_79_21# VPWR 0.017875f
C856 clknet_1_1__leaf_clk hold3/a_285_47# 7.46e-19
C857 _26_/a_634_183# net3 0.002405f
C858 _25_/a_572_47# count[0] 6.77e-19
C859 _27_/a_27_47# _04_ 0.293978f
C860 VPWR clkbuf_1_1__f_clk/a_110_47# 0.330578f
C861 _27_/a_381_47# count[3] 0.01433f
C862 clknet_1_0__leaf_clk _24_/a_475_413# 0.042486f
C863 _21_/a_207_413# _09_ 0.039121f
C864 hold2/a_391_47# _24_/a_193_47# 9.55e-19
C865 _21_/a_297_47# _09_ 0.001026f
C866 net2 clknet_0_clk 0.010995f
C867 _08_ count[3] 0.029923f
C868 net1 clknet_0_clk 0.030715f
C869 hold2/a_285_47# _24_/a_27_47# 0.008609f
C870 _19_/a_561_47# VPWR -3.92e-19
C871 _00_ _25_/a_475_413# 8.78e-20
C872 net3 clkbuf_0_clk/a_110_47# 0.043733f
C873 clknet_1_1__leaf_clk _03_ 0.136016f
C874 _27_/a_891_413# _04_ 0.001417f
C875 _15_/a_297_47# _24_/a_1062_300# 3.11e-19
C876 clknet_1_0__leaf_clk hold1/a_49_47# 6.12e-19
C877 _21_/a_207_413# _10_ 0.001982f
C878 _21_/a_297_47# _10_ 8.27e-19
C879 _15_/a_79_21# net3 4.66e-19
C880 hold2/a_49_47# count[1] 0.001728f
C881 hold1/a_285_47# _24_/a_634_183# 0.010224f
C882 clknet_1_0__leaf_clk count[1] 0.198449f
C883 _26_/a_475_413# VPWR 0.008476f
C884 _24_/a_27_47# clkbuf_1_0__f_clk/a_110_47# 7.58e-19
C885 _26_/a_572_47# VPWR 1.53e-19
C886 _03_ _27_/a_27_47# 6.55e-19
C887 _01_ count[0] 0.010501f
C888 _20_/a_80_21# _06_ 0.002123f
C889 hold3/a_49_47# count[2] 0.037709f
C890 count[0] _24_/a_891_413# 0.037703f
C891 _13_/a_109_297# net4 7.42e-19
C892 _26_/a_891_413# count[0] 0.004702f
C893 count[0] VPWR 1.277962f
C894 hold1/a_285_47# _24_/a_193_47# 0.001481f
C895 net3 _26_/a_475_413# 0.004596f
C896 _09_ VPWR 0.184549f
C897 _27_/a_381_47# _04_ 0.01507f
C898 clknet_1_0__leaf_clk net2 0.005458f
C899 _02_ rst 0.22907f
C900 hold3/a_285_47# _07_ 0.006803f
C901 clknet_1_0__leaf_clk net1 0.15247f
C902 _08_ _04_ 0.035578f
C903 _00_ _04_ 1.52e-19
C904 _10_ VPWR 0.364134f
C905 _21_/a_207_413# clknet_1_1__leaf_clk 2.9e-19
C906 _23_/a_1283_21# _24_/a_1062_300# 0.00786f
C907 _25_/a_1062_300# clknet_1_0__leaf_clk 0.009985f
C908 input1/a_75_212# VPWR 0.093425f
C909 _25_/a_27_47# clknet_0_clk 0.013689f
C910 _03_ _07_ 0.020789f
C911 net3 count[0] 0.689098f
C912 rst net4 1.81e-19
C913 _05_ clknet_0_clk 0.153541f
C914 _15_/a_297_47# clkbuf_0_clk/a_110_47# 9.88e-20
C915 net6 rst 0.072605f
C916 _23_/a_193_47# _24_/a_891_413# 4.13e-20
C917 _23_/a_193_47# VPWR -0.206438f
C918 hold2/a_285_47# _02_ 4.03e-20
C919 _21_/a_207_413# _27_/a_27_47# 2.62e-19
C920 _27_/a_381_47# _03_ 5.54e-21
C921 _25_/a_891_413# count[0] 5.76e-20
C922 _08_ _03_ 2.14e-19
C923 count[3] _26_/a_27_47# 0.1654f
C924 _25_/a_475_413# _02_ 8.56e-19
C925 count[1] _17_/a_209_47# 0.005396f
C926 _23_/a_1462_47# VPWR 2.97e-19
C927 _19_/a_465_47# count[0] 0.001794f
C928 hold2/a_285_47# net4 0.004195f
C929 _02_ clkbuf_1_0__f_clk/a_110_47# 0.007865f
C930 count[1] _14_/a_113_297# 0.019481f
C931 net6 hold2/a_285_47# 3.01e-19
C932 _19_/a_381_47# count[1] 5.56e-19
C933 hold1/a_391_47# count[0] 0.008124f
C934 _26_/a_193_47# clkbuf_0_clk/a_110_47# 1.32e-19
C935 clknet_1_1__leaf_clk _26_/a_891_413# 7.78e-19
C936 _24_/a_572_47# VPWR 8.18e-21
C937 _27_/a_193_47# _27_/a_634_183# -0.001855f
C938 _25_/a_475_413# net6 7.49e-19
C939 clknet_1_1__leaf_clk VPWR 0.337343f
C940 count[2] _19_/a_79_21# 0.004038f
C941 net2 _23_/a_448_47# 0.006776f
C942 _25_/a_193_47# _24_/a_891_413# 5.66e-20
C943 _26_/a_634_183# count[2] 0.005019f
C944 _25_/a_27_47# clknet_1_0__leaf_clk 0.435702f
C945 net1 _23_/a_448_47# 0.016613f
C946 _05_ clknet_1_0__leaf_clk 9.24e-20
C947 _25_/a_193_47# VPWR 0.008812f
C948 _26_/a_193_47# clkbuf_1_1__f_clk/a_110_47# 1.24e-20
C949 net4 clkbuf_1_0__f_clk/a_110_47# 1.49e-19
C950 net6 clkbuf_1_0__f_clk/a_110_47# 3.99e-19
C951 _27_/a_568_413# clknet_0_clk 6.57e-19
C952 clkbuf_0_clk/a_110_47# count[2] 0.00706f
C953 clknet_1_0__leaf_clk _17_/a_80_21# 3.56e-20
C954 _27_/a_27_47# VPWR -0.180488f
C955 _21_/a_27_413# count[1] 8.43e-19
C956 _15_/a_297_47# count[0] 0.018792f
C957 _21_/a_27_413# _27_/a_193_47# 6.84e-19
C958 _26_/a_27_47# _04_ 6.25e-19
C959 clkbuf_1_1__f_clk/a_110_47# count[2] 0.003811f
C960 _21_/a_297_47# _08_ 9.16e-19
C961 _21_/a_207_413# _08_ 0.005849f
C962 net3 _25_/a_193_47# 7.42e-20
C963 _26_/a_475_413# _26_/a_193_47# -0.003877f
C964 _27_/a_891_413# VPWR 0.0122f
C965 _19_/a_561_47# count[2] 5.25e-19
C966 _22_/a_75_212# clk 6.79e-21
C967 _10_ _20_/a_209_47# 2.14e-19
C968 hold4/a_49_47# _24_/a_27_47# 2.05e-19
C969 _26_/a_891_413# _07_ 0.01623f
C970 _16_/a_199_47# _20_/a_80_21# 1.16e-20
C971 _26_/a_193_47# count[0] 0.032265f
C972 count[3] _27_/a_475_413# 0.031904f
C973 _26_/a_475_413# count[2] 0.003143f
C974 _06_ hold3/a_391_47# 0.001715f
C975 _17_/a_209_297# count[0] 0.004736f
C976 _07_ VPWR 0.210351f
C977 count[1] _25_/a_381_47# 8.74e-20
C978 rst clknet_0_clk 0.267149f
C979 _03_ _26_/a_27_47# 0.082513f
C980 _26_/a_381_47# count[3] 0.010793f
C981 _23_/a_1283_21# count[0] 6.93e-19
C982 clknet_1_0__leaf_clk _24_/a_975_413# 0.00206f
C983 _01_ _24_/a_27_47# 1.21e-20
C984 _27_/a_381_47# VPWR -0.001652f
C985 count[0] count[2] 0.527532f
C986 _00_ _24_/a_891_413# 1.98e-19
C987 _27_/a_1062_300# _10_ 0.024329f
C988 _08_ VPWR 0.340963f
C989 count[1] _24_/a_475_413# 0.027724f
C990 _00_ VPWR 0.175098f
C991 _25_/a_634_183# _24_/a_1062_300# 5.17e-19
C992 _09_ count[2] 0.004003f
C993 net6 _03_ 0.001737f
C994 net3 _07_ 7.3e-19
C995 _05_ _14_/a_113_297# 0.005084f
C996 _24_/a_27_47# VPWR -0.070711f
C997 _16_/a_113_297# count[1] 0.002581f
C998 _17_/a_80_21# _14_/a_113_297# 6.73e-20
C999 count[1] hold1/a_49_47# 0.005636f
C1000 _10_ count[2] 0.002655f
C1001 _25_/a_475_413# clknet_0_clk 3.26e-19
C1002 _17_/a_303_47# count[0] 1.78e-19
C1003 count[3] clknet_0_clk 0.024143f
C1004 _15_/a_297_47# _25_/a_193_47# 6.24e-21
C1005 _23_/a_543_47# count[0] 2.45e-20
C1006 hold2/a_49_47# rst 2.95e-21
C1007 _08_ net3 4.12e-20
C1008 _27_/a_475_413# _04_ 0.040621f
C1009 _23_/a_27_47# _23_/a_761_289# -6.54e-19
C1010 clknet_1_0__leaf_clk rst 0.001558f
C1011 _10_ _27_/a_975_413# 0.00107f
C1012 clknet_0_clk clkbuf_1_0__f_clk/a_110_47# 0.00666f
C1013 count[0] _24_/a_1020_47# 5.96e-19
C1014 net3 _24_/a_27_47# 7.61e-19
C1015 _26_/a_381_47# _04_ 3.1e-22
C1016 _23_/a_1108_47# _24_/a_193_47# 2.04e-20
C1017 clknet_1_1__leaf_clk _26_/a_193_47# 0.286269f
C1018 _25_/a_1062_300# _24_/a_475_413# 0.007354f
C1019 _27_/a_1062_300# clknet_1_1__leaf_clk 1.81e-19
C1020 _25_/a_891_413# _24_/a_27_47# 0.011052f
C1021 net5 hold3/a_391_47# 0.006599f
C1022 hold4/a_49_47# net4 0.001457f
C1023 _23_/a_193_47# _23_/a_543_47# -0.012086f
C1024 hold2/a_285_47# clknet_1_0__leaf_clk 0.014157f
C1025 net6 hold4/a_49_47# 6.52e-19
C1026 _03_ _27_/a_475_413# 8.39e-21
C1027 _25_/a_634_183# clkbuf_0_clk/a_110_47# 1.57e-19
C1028 _27_/a_27_47# _26_/a_193_47# 7.18e-19
C1029 clknet_1_1__leaf_clk count[2] 0.064816f
C1030 _26_/a_1062_300# hold3/a_391_47# 0.010284f
C1031 _25_/a_1062_300# count[1] 0.061046f
C1032 _25_/a_475_413# clknet_1_0__leaf_clk 0.044202f
C1033 hold1/a_391_47# _24_/a_27_47# 9.29e-19
C1034 _04_ clknet_0_clk 0.197756f
C1035 _03_ _26_/a_381_47# 0.020813f
C1036 _19_/a_297_297# _19_/a_79_21# -6.12e-20
C1037 _25_/a_27_47# _25_/a_381_47# -0.004383f
C1038 net5 _06_ 0.160451f
C1039 _05_ _25_/a_381_47# 5.36e-19
C1040 hold1/a_285_47# hold2/a_391_47# 3.65e-19
C1041 count[0] _26_/a_568_413# 0.001641f
C1042 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# 0.05153f
C1043 net1 net2 0.021363f
C1044 _02_ VPWR 0.468554f
C1045 _19_/a_297_297# clkbuf_0_clk/a_110_47# 3.72e-19
C1046 _26_/a_27_47# VPWR -0.0604f
C1047 _27_/a_27_47# count[2] 0.007689f
C1048 _26_/a_1062_300# _06_ 0.009941f
C1049 n_rst clknet_1_0__leaf_clk 0.005322f
C1050 _27_/a_1020_47# count[3] 5.98e-19
C1051 _08_ _20_/a_209_47# 9.07e-19
C1052 _18_/a_109_297# _06_ 9.49e-19
C1053 _01_ net4 0.00339f
C1054 _23_/a_448_47# rst 9.03e-20
C1055 net6 _01_ 0.002444f
C1056 _05_ _24_/a_475_413# 1.19e-20
C1057 net4 _24_/a_891_413# 6.49e-20
C1058 count[0] _24_/a_634_183# 0.003661f
C1059 net6 _24_/a_891_413# 0.035861f
C1060 _03_ clknet_0_clk 5.15e-19
C1061 _07_ _26_/a_193_47# 5.3e-19
C1062 net4 VPWR 0.046103f
C1063 _17_/a_80_21# _24_/a_475_413# 1.63e-21
C1064 net6 VPWR 0.101083f
C1065 _07_ _17_/a_209_297# 0.002255f
C1066 net3 _26_/a_27_47# 2.72e-19
C1067 hold4/a_391_47# _24_/a_27_47# 0.001156f
C1068 _19_/a_381_47# rst 6.59e-19
C1069 _05_ hold1/a_49_47# 1.65e-19
C1070 _20_/a_80_21# clkbuf_0_clk/a_110_47# 4.51e-20
C1071 net3 _02_ 2.14e-19
C1072 _23_/a_761_289# count[0] 6.67e-20
C1073 _21_/a_207_413# _27_/a_475_413# 5.02e-19
C1074 _25_/a_27_47# count[1] 0.003199f
C1075 _17_/a_80_21# hold1/a_49_47# 2.07e-20
C1076 _05_ count[1] 0.008701f
C1077 _08_ _26_/a_193_47# 7.1e-19
C1078 _25_/a_634_183# count[0] 0.007555f
C1079 _24_/a_193_47# count[0] 0.004522f
C1080 _07_ count[2] 0.211454f
C1081 _20_/a_80_21# clkbuf_1_1__f_clk/a_110_47# 2.51e-20
C1082 _23_/a_651_413# VPWR -0.009331f
C1083 _25_/a_891_413# _02_ 3.43e-19
C1084 _08_ _17_/a_209_297# 9.88e-20
C1085 net3 net4 0.078403f
C1086 _17_/a_80_21# count[1] 0.111425f
C1087 _16_/a_199_47# _06_ -2.22e-34
C1088 net6 net3 6.7e-19
C1089 _10_ _23_/a_761_289# 8.74e-20
C1090 _27_/a_381_47# count[2] 1.67e-21
C1091 _15_/a_382_297# count[0] 9.21e-19
C1092 _08_ count[2] 0.074858f
C1093 _00_ _23_/a_1283_21# 3.53e-19
C1094 hold1/a_391_47# _02_ 3.39e-19
C1095 _19_/a_297_297# count[0] 0.011363f
C1096 clknet_1_1__leaf_clk _26_/a_568_413# 1.34e-19
C1097 hold1/a_391_47# _26_/a_27_47# 3.19e-21
C1098 _25_/a_27_47# net1 1.57e-19
C1099 _25_/a_891_413# net6 3.1e-21
C1100 _23_/a_1270_413# count[0] 1.43e-20
C1101 _23_/a_1283_21# _24_/a_27_47# 6.82e-20
C1102 count[3] _27_/a_634_183# 0.01585f
C1103 n_rst _23_/a_448_47# 6.64e-20
C1104 _23_/a_193_47# _23_/a_761_289# -0.00122f
C1105 _21_/a_207_413# clknet_0_clk 0.017368f
C1106 _21_/a_297_47# clknet_0_clk 9.15e-19
C1107 _25_/a_572_47# clknet_0_clk 9.65e-20
C1108 _23_/a_193_47# _24_/a_193_47# 2.49e-20
C1109 _27_/a_475_413# VPWR 0.003428f
C1110 hold1/a_391_47# net4 0.001685f
C1111 _26_/a_1062_300# net5 4.58e-19
C1112 net6 hold1/a_391_47# 4.47e-20
C1113 _18_/a_109_297# net5 0.002068f
C1114 _24_/a_381_47# VPWR -0.002848f
C1115 _20_/a_80_21# count[0] 0.024666f
C1116 _26_/a_381_47# VPWR 0.001495f
C1117 _00_ _23_/a_543_47# 0.01009f
C1118 _21_/a_27_413# count[3] 1.49e-19
C1119 _25_/a_193_47# _24_/a_634_183# 8.84e-20
C1120 hold3/a_49_47# _06_ 4.9e-19
C1121 _09_ _20_/a_80_21# 8.26e-19
C1122 _20_/a_303_47# VPWR -4.38e-19
C1123 _27_/a_572_47# _08_ 5.22e-19
C1124 count[1] _24_/a_975_413# 4.04e-19
C1125 _13_/a_109_297# count[1] 0.001581f
C1126 _24_/a_193_47# _24_/a_572_47# -9.97e-19
C1127 _01_ clknet_0_clk 6.36e-20
C1128 _10_ _20_/a_80_21# 1.07e-19
C1129 _15_/a_297_47# net4 1.79e-19
C1130 net6 _15_/a_297_47# 0.013591f
C1131 _22_/a_75_212# _19_/a_79_21# 2.28e-20
C1132 _25_/a_634_183# _25_/a_193_47# -0.001855f
C1133 _24_/a_891_413# clknet_0_clk 1.22e-20
C1134 _25_/a_193_47# _24_/a_193_47# 3.47e-20
C1135 _04_ _27_/a_634_183# 0.023269f
C1136 hold4/a_391_47# net4 0.003533f
C1137 _26_/a_27_47# _26_/a_193_47# -0.096811f
C1138 VPWR clknet_0_clk 1.27397f
C1139 net6 hold4/a_391_47# 0.001565f
C1140 clknet_1_0__leaf_clk hold4/a_49_47# 2.21e-19
C1141 _25_/a_27_47# _05_ 2.88e-20
C1142 hold1/a_49_47# rst 0.007504f
C1143 clknet_1_1__leaf_clk _19_/a_297_297# 5.09e-19
C1144 _17_/a_209_297# _26_/a_27_47# 6.57e-19
C1145 _25_/a_568_413# count[0] 8.25e-19
C1146 count[1] rst 0.01255f
C1147 _21_/a_27_413# _04_ 0.002527f
C1148 _02_ _23_/a_1283_21# 0.004039f
C1149 net6 _26_/a_193_47# 4.55e-21
C1150 _26_/a_27_47# count[2] 0.048143f
C1151 _25_/a_381_47# clkbuf_1_0__f_clk/a_110_47# 9.78e-19
C1152 net3 clknet_0_clk 0.115144f
C1153 _02_ count[2] 0.002895f
C1154 hold2/a_49_47# _01_ 0.049789f
C1155 _03_ _27_/a_634_183# 1.81e-21
C1156 clknet_1_1__leaf_clk _20_/a_80_21# 0.015056f
C1157 _16_/a_113_297# count[3] 2.16e-20
C1158 hold2/a_49_47# VPWR 0.066914f
C1159 _24_/a_475_413# clkbuf_1_0__f_clk/a_110_47# 8.21e-19
C1160 clknet_1_0__leaf_clk _24_/a_891_413# 0.036555f
C1161 _25_/a_475_413# hold1/a_49_47# 2.73e-20
C1162 net6 _23_/a_1283_21# 1.05e-20
C1163 net4 count[2] 4.84e-20
C1164 net6 count[2] 2.07e-20
C1165 _00_ _24_/a_634_183# 1.58e-20
C1166 net2 rst 8.61e-20
C1167 net1 rst 1.03e-19
C1168 hold2/a_285_47# count[1] 0.008831f
C1169 clknet_1_0__leaf_clk VPWR 1.562421f
C1170 hold3/a_49_47# net5 6.42e-19
C1171 _24_/a_27_47# _24_/a_634_183# -0.004305f
C1172 _25_/a_475_413# count[1] 2.98e-19
C1173 count[3] count[1] 0.169548f
C1174 _23_/a_1108_47# clk 1.14e-19
C1175 _23_/a_27_47# clk 0.001735f
C1176 _14_/a_199_47# clknet_0_clk 4.23e-20
C1177 count[3] _27_/a_193_47# 0.028087f
C1178 hold1/a_49_47# clkbuf_1_0__f_clk/a_110_47# 5.56e-22
C1179 _27_/a_27_47# _20_/a_80_21# 1.55e-19
C1180 _00_ _23_/a_761_289# 0.013767f
C1181 count[1] clkbuf_1_0__f_clk/a_110_47# 0.036588f
C1182 hold2/a_49_47# net3 3.83e-19
C1183 _22_/a_75_212# count[0] 1.04e-19
C1184 _07_ _19_/a_297_297# 2.03e-19
C1185 _00_ _25_/a_634_183# 6.47e-21
C1186 _00_ _24_/a_193_47# 0.001502f
C1187 _27_/a_1020_47# VPWR -4.43e-19
C1188 net3 clknet_1_0__leaf_clk 6.73e-20
C1189 _24_/a_193_47# _24_/a_27_47# -0.158901f
C1190 _25_/a_634_183# _24_/a_27_47# 8.67e-20
C1191 _05_ _13_/a_109_297# 2.89e-19
C1192 count[0] _24_/a_568_413# 1.67e-19
C1193 count[3] net2 4.56e-21
C1194 clk clkbuf_0_clk/a_110_47# 0.004735f
C1195 net6 _24_/a_1020_47# 0.001851f
C1196 _21_/a_207_413# _27_/a_634_183# 0.006947f
C1197 _08_ _19_/a_297_297# 0.002087f
C1198 _10_ _22_/a_75_212# 0.054952f
C1199 _26_/a_381_47# _26_/a_193_47# -0.004383f
C1200 _25_/a_891_413# clknet_1_0__leaf_clk 0.011723f
C1201 _00_ _23_/a_1270_413# 1.62e-19
C1202 n_rst net2 3.45e-19
C1203 count[1] _04_ 5.23e-20
C1204 count[0] hold3/a_391_47# 6.95e-19
C1205 n_rst net1 0.003766f
C1206 _23_/a_1217_47# clknet_0_clk 3.45e-19
C1207 _27_/a_193_47# _04_ 0.178479f
C1208 _25_/a_1062_300# clkbuf_1_0__f_clk/a_110_47# 0.034938f
C1209 hold3/a_285_47# _16_/a_113_297# 3.51e-19
C1210 hold1/a_391_47# clknet_1_0__leaf_clk 5.65e-20
C1211 _25_/a_27_47# rst 4.74e-21
C1212 _23_/a_448_47# VPWR -0.002712f
C1213 _26_/a_381_47# count[2] 8.34e-21
C1214 _05_ rst 0.124131f
C1215 _01_ _14_/a_113_297# 0.001095f
C1216 _08_ _20_/a_80_21# 0.025603f
C1217 VPWR _17_/a_209_47# -0.001019f
C1218 _20_/a_303_47# count[2] 0.005211f
C1219 hold3/a_285_47# count[1] 1.17e-19
C1220 _03_ _16_/a_113_297# 0.009398f
C1221 count[0] _06_ 0.030764f
C1222 _26_/a_891_413# _14_/a_113_297# 7.41e-21
C1223 VPWR _14_/a_113_297# 0.070686f
C1224 _19_/a_381_47# VPWR 0.00185f
C1225 _09_ _06_ 9.87e-21
C1226 VPWR _27_/a_634_183# 6.71e-19
C1227 _03_ count[1] 0.384241f
C1228 net3 _17_/a_209_47# 0.001251f
C1229 _03_ _27_/a_193_47# 2.01e-19
C1230 hold2/a_391_47# count[0] 3.86e-19
C1231 _23_/a_1283_21# clknet_0_clk 0.019248f
C1232 count[0] clk 7.27e-20
C1233 clknet_0_clk count[2] 0.010709f
C1234 _25_/a_475_413# _25_/a_27_47# -0.01416f
C1235 hold2/a_49_47# hold4/a_391_47# 3.2e-19
C1236 net4 _24_/a_634_183# 3.11e-19
C1237 _25_/a_475_413# _05_ 2.84e-22
C1238 net6 _24_/a_634_183# 0.02234f
C1239 _05_ count[3] 0.003688f
C1240 clknet_1_0__leaf_clk hold4/a_391_47# 0.013378f
C1241 net3 _14_/a_113_297# 0.006211f
C1242 _02_ _24_/a_193_47# 3.91e-20
C1243 _25_/a_634_183# _02_ 6.07e-19
C1244 count[3] _17_/a_80_21# 1.23e-19
C1245 _22_/a_75_212# _27_/a_27_47# 5.59e-19
C1246 _21_/a_27_413# VPWR -4.77e-19
C1247 _25_/a_27_47# clkbuf_1_0__f_clk/a_110_47# 0.013722f
C1248 _05_ clkbuf_1_0__f_clk/a_110_47# 1.67e-19
C1249 _10_ clk 1.65e-19
C1250 _00_ _25_/a_568_413# 2.73e-20
C1251 input1/a_75_212# clk 0.00167f
C1252 _23_/a_543_47# clknet_0_clk 0.001715f
C1253 _25_/a_891_413# _14_/a_113_297# 5.94e-21
C1254 _15_/a_382_297# _02_ 3.37e-19
C1255 VPWR VGND 0.22244p
C1256 _00_ VGND 0.346385f
C1257 net1 VGND 0.587444f
C1258 _13_/a_109_297# VGND -5.49e-19
C1259 _14_/a_199_47# VGND 0.001592f
C1260 _14_/a_113_297# VGND 0.047168f
C1261 net6 VGND 1.145445f
C1262 _05_ VGND 0.198598f
C1263 _15_/a_297_47# VGND 0.037191f
C1264 _15_/a_382_297# VGND -4.43e-19
C1265 _15_/a_79_21# VGND 0.162256f
C1266 clkbuf_1_1__f_clk/a_110_47# VGND 1.987437f
C1267 _06_ VGND 0.171859f
C1268 net5 VGND 0.30965f
C1269 _16_/a_199_47# VGND -2.37e-19
C1270 _16_/a_113_297# VGND 0.045032f
C1271 _23__2/LO VGND 0.267239f
C1272 _07_ VGND 0.412929f
C1273 _17_/a_303_47# VGND 0.001601f
C1274 _17_/a_209_47# VGND 0.004632f
C1275 _17_/a_209_297# VGND 0.0166f
C1276 _17_/a_80_21# VGND 0.243138f
C1277 hold4/a_391_47# VGND 0.148028f
C1278 hold4/a_285_47# VGND 0.347943f
C1279 hold4/a_49_47# VGND 0.38987f
C1280 _18_/a_109_297# VGND 0.002775f
C1281 hold3/a_391_47# VGND 0.150121f
C1282 hold3/a_285_47# VGND 0.346013f
C1283 hold3/a_49_47# VGND 0.357301f
C1284 _08_ VGND 0.391403f
C1285 count[2] VGND 2.348828f
C1286 _19_/a_561_47# VGND -5.95e-19
C1287 _19_/a_465_47# VGND -8.41e-19
C1288 _19_/a_381_47# VGND -4.51e-19
C1289 _19_/a_297_297# VGND 0.032008f
C1290 _19_/a_79_21# VGND 0.144337f
C1291 _01_ VGND 0.345625f
C1292 hold2/a_391_47# VGND 0.135243f
C1293 hold2/a_285_47# VGND 0.308755f
C1294 hold2/a_49_47# VGND 0.354323f
C1295 net3 VGND 0.931803f
C1296 hold1/a_391_47# VGND 0.180268f
C1297 hold1/a_285_47# VGND 0.363191f
C1298 hold1/a_49_47# VGND 0.311005f
C1299 clknet_1_0__leaf_clk VGND 1.724413f
C1300 clknet_0_clk VGND 3.041779f
C1301 clkbuf_1_0__f_clk/a_110_47# VGND 1.980781f
C1302 n_rst VGND 0.554047f
C1303 input1/a_75_212# VGND 0.278906f
C1304 _09_ VGND 0.206056f
C1305 _20_/a_303_47# VGND 1.18e-19
C1306 _20_/a_209_47# VGND -1.41e-19
C1307 _20_/a_209_297# VGND 0.005621f
C1308 _20_/a_80_21# VGND 0.224181f
C1309 _21_/a_297_47# VGND 3.54e-19
C1310 _21_/a_207_413# VGND 0.161646f
C1311 _21_/a_27_413# VGND 0.20938f
C1312 _04_ VGND 0.238975f
C1313 _10_ VGND 0.760316f
C1314 _22_/a_75_212# VGND 0.26029f
C1315 rst VGND 0.812577f
C1316 net2 VGND 0.721089f
C1317 _23_/a_1462_47# VGND 2.59e-19
C1318 _23_/a_1217_47# VGND 1.43e-19
C1319 _23_/a_805_47# VGND 0.002795f
C1320 _23_/a_639_47# VGND 0.004739f
C1321 _23_/a_1270_413# VGND 7.79e-20
C1322 _23_/a_651_413# VGND 0.014975f
C1323 _23_/a_448_47# VGND 0.018341f
C1324 _23_/a_1108_47# VGND 0.157514f
C1325 _23_/a_1283_21# VGND 0.31902f
C1326 _23_/a_543_47# VGND 0.184013f
C1327 _23_/a_761_289# VGND 0.140587f
C1328 _23_/a_193_47# VGND 0.323115f
C1329 _23_/a_27_47# VGND 0.56521f
C1330 count[0] VGND 2.544707f
C1331 net4 VGND 0.327057f
C1332 _24_/a_1020_47# VGND -2.22e-19
C1333 _24_/a_572_47# VGND 0.001226f
C1334 _24_/a_975_413# VGND -2.21e-19
C1335 _24_/a_568_413# VGND 0.002046f
C1336 _24_/a_381_47# VGND 0.014193f
C1337 _24_/a_891_413# VGND 0.149083f
C1338 _24_/a_1062_300# VGND 0.522403f
C1339 _24_/a_475_413# VGND 0.158032f
C1340 _24_/a_634_183# VGND 0.174418f
C1341 _24_/a_193_47# VGND 0.075569f
C1342 _24_/a_27_47# VGND 0.501827f
C1343 clk VGND 1.629049f
C1344 clkbuf_0_clk/a_110_47# VGND 1.77177f
C1345 count[1] VGND 3.160929f
C1346 _02_ VGND 0.365319f
C1347 _25_/a_1020_47# VGND 0.002448f
C1348 _25_/a_572_47# VGND 2.7e-19
C1349 _25_/a_975_413# VGND 0.002645f
C1350 _25_/a_568_413# VGND 3.3e-19
C1351 _25_/a_381_47# VGND 0.018191f
C1352 _25_/a_891_413# VGND 0.197662f
C1353 _25_/a_1062_300# VGND 0.580156f
C1354 _25_/a_475_413# VGND 0.140942f
C1355 _25_/a_634_183# VGND 0.154405f
C1356 _25_/a_193_47# VGND 0.294393f
C1357 _25_/a_27_47# VGND 0.485801f
C1358 _03_ VGND 0.567601f
C1359 _26_/a_1020_47# VGND 0.002315f
C1360 _26_/a_572_47# VGND 1.85e-19
C1361 _26_/a_975_413# VGND 0.002012f
C1362 _26_/a_568_413# VGND 1.99e-19
C1363 _26_/a_381_47# VGND 0.017982f
C1364 _26_/a_891_413# VGND 0.180222f
C1365 _26_/a_1062_300# VGND 0.594146f
C1366 _26_/a_475_413# VGND 0.143042f
C1367 _26_/a_634_183# VGND 0.159981f
C1368 _26_/a_193_47# VGND 0.318152f
C1369 _26_/a_27_47# VGND 0.495614f
C1370 count[3] VGND 1.231933f
C1371 clknet_1_1__leaf_clk VGND 0.863186f
C1372 _27_/a_1020_47# VGND 0.002047f
C1373 _27_/a_572_47# VGND 2.56e-19
C1374 _27_/a_975_413# VGND 3.42e-19
C1375 _27_/a_568_413# VGND 2.48e-19
C1376 _27_/a_381_47# VGND 0.017857f
C1377 _27_/a_891_413# VGND 0.191179f
C1378 _27_/a_1062_300# VGND 0.645405f
C1379 _27_/a_475_413# VGND 0.147025f
C1380 _27_/a_634_183# VGND 0.165334f
C1381 _27_/a_193_47# VGND 0.292484f
C1382 _27_/a_27_47# VGND 0.494967f
.ends

